VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_greycode_top
  CLASS BLOCK ;
  FOREIGN tt_um_greycode_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 679.880 BY 220.320 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 219.150 158.850 220.320 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 162.230 219.320 162.530 220.320 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 216.740 155.170 220.320 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 218.780 151.490 220.320 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 216.740 147.810 220.320 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 216.740 144.130 220.320 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 218.780 140.450 220.320 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 214.020 136.770 220.320 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 218.780 133.090 220.320 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 214.020 129.410 220.320 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 215.380 125.730 220.320 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 218.100 122.050 220.320 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 216.740 118.370 220.320 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 215.380 114.690 220.320 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 214.020 111.010 220.320 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 214.020 107.330 220.320 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 218.780 103.650 220.320 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 218.780 99.970 220.320 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 218.780 96.290 220.320 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 211.980 33.730 220.320 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 211.980 30.050 220.320 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 214.700 26.370 220.320 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 216.060 22.690 220.320 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 214.700 19.010 220.320 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 218.780 15.330 220.320 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 211.980 11.650 220.320 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 218.780 7.970 220.320 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 218.780 63.170 220.320 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 218.780 59.490 220.320 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 218.780 55.810 220.320 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 218.780 52.130 220.320 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 214.700 48.450 220.320 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 214.700 44.770 220.320 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 218.780 41.090 220.320 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 218.100 37.410 220.320 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 218.100 92.610 220.320 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 218.100 88.930 220.320 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 218.780 85.250 220.320 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 218.780 81.570 220.320 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 218.780 77.890 220.320 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 218.780 74.210 220.320 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 218.780 70.530 220.320 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 218.100 66.850 220.320 ;
    END
  END uo_out[7]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 5.200 22.640 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 5.200 176.240 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 5.200 329.840 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 5.200 483.440 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 5.200 637.040 215.120 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 5.200 99.440 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 5.200 253.040 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 5.200 406.640 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 5.200 560.240 215.120 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 213.465 674.550 215.070 ;
        RECT 5.330 208.025 674.550 210.855 ;
        RECT 5.330 202.585 674.550 205.415 ;
        RECT 5.330 197.145 674.550 199.975 ;
        RECT 5.330 191.705 674.550 194.535 ;
        RECT 5.330 186.265 674.550 189.095 ;
        RECT 5.330 180.825 674.550 183.655 ;
        RECT 5.330 175.385 674.550 178.215 ;
        RECT 5.330 169.945 674.550 172.775 ;
        RECT 5.330 164.505 674.550 167.335 ;
        RECT 5.330 159.065 674.550 161.895 ;
        RECT 5.330 153.625 674.550 156.455 ;
        RECT 5.330 148.185 674.550 151.015 ;
        RECT 5.330 142.745 674.550 145.575 ;
        RECT 5.330 137.305 674.550 140.135 ;
        RECT 5.330 131.865 674.550 134.695 ;
        RECT 5.330 126.425 674.550 129.255 ;
        RECT 5.330 120.985 674.550 123.815 ;
        RECT 5.330 115.545 674.550 118.375 ;
        RECT 5.330 110.105 674.550 112.935 ;
        RECT 5.330 104.665 674.550 107.495 ;
        RECT 5.330 99.225 674.550 102.055 ;
        RECT 5.330 93.785 674.550 96.615 ;
        RECT 5.330 88.345 674.550 91.175 ;
        RECT 5.330 82.905 674.550 85.735 ;
        RECT 5.330 77.465 674.550 80.295 ;
        RECT 5.330 72.025 674.550 74.855 ;
        RECT 5.330 66.585 674.550 69.415 ;
        RECT 5.330 61.145 674.550 63.975 ;
        RECT 5.330 55.705 674.550 58.535 ;
        RECT 5.330 50.265 674.550 53.095 ;
        RECT 5.330 44.825 674.550 47.655 ;
        RECT 5.330 39.385 674.550 42.215 ;
        RECT 5.330 33.945 674.550 36.775 ;
        RECT 5.330 28.505 674.550 31.335 ;
        RECT 5.330 23.065 674.550 25.895 ;
        RECT 5.330 17.625 674.550 20.455 ;
        RECT 5.330 12.185 674.550 15.015 ;
        RECT 5.330 6.745 674.550 9.575 ;
      LAYER li1 ;
        RECT 5.520 5.355 674.360 214.965 ;
      LAYER met1 ;
        RECT 5.520 5.200 674.360 217.900 ;
      LAYER met2 ;
        RECT 9.300 5.255 671.040 218.805 ;
      LAYER met3 ;
        RECT 7.630 5.275 637.030 218.785 ;
      LAYER met4 ;
        RECT 8.370 218.380 10.950 219.450 ;
        RECT 7.655 211.580 10.950 218.380 ;
        RECT 12.050 218.380 14.630 219.450 ;
        RECT 15.730 218.380 18.310 219.450 ;
        RECT 12.050 214.300 18.310 218.380 ;
        RECT 19.410 215.660 21.990 219.450 ;
        RECT 23.090 215.660 25.670 219.450 ;
        RECT 19.410 215.520 25.670 215.660 ;
        RECT 19.410 214.300 20.640 215.520 ;
        RECT 12.050 211.580 20.640 214.300 ;
        RECT 7.655 193.295 20.640 211.580 ;
        RECT 23.040 214.300 25.670 215.520 ;
        RECT 26.770 214.300 29.350 219.450 ;
        RECT 23.040 211.580 29.350 214.300 ;
        RECT 30.450 211.580 33.030 219.450 ;
        RECT 34.130 217.700 36.710 219.450 ;
        RECT 37.810 218.380 40.390 219.450 ;
        RECT 41.490 218.380 44.070 219.450 ;
        RECT 37.810 217.700 44.070 218.380 ;
        RECT 34.130 214.300 44.070 217.700 ;
        RECT 45.170 214.300 47.750 219.450 ;
        RECT 48.850 218.380 51.430 219.450 ;
        RECT 52.530 218.380 55.110 219.450 ;
        RECT 56.210 218.380 58.790 219.450 ;
        RECT 59.890 218.380 62.470 219.450 ;
        RECT 63.570 218.380 66.150 219.450 ;
        RECT 48.850 217.700 66.150 218.380 ;
        RECT 67.250 218.380 69.830 219.450 ;
        RECT 70.930 218.380 73.510 219.450 ;
        RECT 74.610 218.380 77.190 219.450 ;
        RECT 78.290 218.380 80.870 219.450 ;
        RECT 81.970 218.380 84.550 219.450 ;
        RECT 85.650 218.380 88.230 219.450 ;
        RECT 67.250 217.700 88.230 218.380 ;
        RECT 89.330 217.700 91.910 219.450 ;
        RECT 93.010 218.380 95.590 219.450 ;
        RECT 96.690 218.380 99.270 219.450 ;
        RECT 100.370 218.380 102.950 219.450 ;
        RECT 104.050 218.380 106.630 219.450 ;
        RECT 93.010 217.700 106.630 218.380 ;
        RECT 48.850 215.520 106.630 217.700 ;
        RECT 48.850 214.300 97.440 215.520 ;
        RECT 34.130 211.580 97.440 214.300 ;
        RECT 23.040 193.295 97.440 211.580 ;
        RECT 99.840 213.620 106.630 215.520 ;
        RECT 107.730 213.620 110.310 219.450 ;
        RECT 111.410 214.980 113.990 219.450 ;
        RECT 115.090 216.340 117.670 219.450 ;
        RECT 118.770 217.700 121.350 219.450 ;
        RECT 122.450 217.700 125.030 219.450 ;
        RECT 118.770 216.340 125.030 217.700 ;
        RECT 115.090 214.980 125.030 216.340 ;
        RECT 126.130 214.980 128.710 219.450 ;
        RECT 111.410 213.620 128.710 214.980 ;
        RECT 129.810 218.380 132.390 219.450 ;
        RECT 133.490 218.380 136.070 219.450 ;
        RECT 129.810 213.620 136.070 218.380 ;
        RECT 137.170 218.380 139.750 219.450 ;
        RECT 140.850 218.380 143.430 219.450 ;
        RECT 137.170 216.340 143.430 218.380 ;
        RECT 144.530 216.340 147.110 219.450 ;
        RECT 148.210 218.380 150.790 219.450 ;
        RECT 151.890 218.380 154.470 219.450 ;
        RECT 148.210 216.340 154.470 218.380 ;
        RECT 155.570 218.750 158.150 219.450 ;
        RECT 159.250 218.750 159.785 219.450 ;
        RECT 155.570 216.340 159.785 218.750 ;
        RECT 137.170 213.620 159.785 216.340 ;
        RECT 99.840 193.295 159.785 213.620 ;
  END
END tt_um_greycode_top
END LIBRARY

