module user_project_wrapper (user_clock2,
    vccd1,
    vccd2,
    vdda1,
    vdda2,
    vssa1,
    vssa2,
    vssd1,
    vssd2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    analog_io,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input vccd1;
 input vccd2;
 input vdda1;
 input vdda2;
 input vssa1;
 input vssa2;
 input vssd1;
 input vssd2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 inout [28:0] analog_io;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire \tt_top1.io_oeb[0] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.clk ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ena ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[10] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[11] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[12] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[13] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[14] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[15] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[16] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[17] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[1] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[2] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[3] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[4] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[5] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[6] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[7] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[8] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[9] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.k_zero ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[0] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[10] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[11] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[12] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[13] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[14] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[15] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[16] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[17] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[18] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[19] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[1] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[20] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[21] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[22] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[23] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[2] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[3] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[4] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[5] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[6] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[7] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[8] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[9] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.clk ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ena ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[10] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[11] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[12] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[13] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[14] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[15] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[16] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[17] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[1] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[2] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[3] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[4] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[5] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[6] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[7] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[8] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[9] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.k_zero ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[0] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[10] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[11] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[12] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[13] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[14] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[15] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[16] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[17] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[18] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[19] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[1] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[20] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[21] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[22] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[23] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[2] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[3] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[4] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[5] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[6] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[7] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[8] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[9] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.clk ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ena ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[10] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[11] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[12] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[13] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[14] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[15] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[16] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[17] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[1] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[2] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[3] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[4] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[5] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[6] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[7] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[8] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[9] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.k_zero ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[0] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[10] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[11] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[12] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[13] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[14] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[15] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[16] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[17] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[18] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[19] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[1] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[20] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[21] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[22] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[23] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[2] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[3] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[4] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[5] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[6] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[7] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[8] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[9] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.clk ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ena ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[10] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[11] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[12] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[13] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[14] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[15] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[16] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[17] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[1] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[2] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[3] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[4] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[5] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[6] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[7] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[8] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[9] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.k_zero ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[0] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[10] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[11] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[12] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[13] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[14] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[15] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[16] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[17] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[18] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[19] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[1] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[20] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[21] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[22] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[23] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[2] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[3] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[4] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[5] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[6] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[7] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[8] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[9] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.clk ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ena ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[10] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[11] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[12] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[13] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[14] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[15] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[16] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[17] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[1] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[2] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[3] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[4] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[5] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[6] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[7] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[8] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[9] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.k_zero ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[0] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[10] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[11] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[12] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[13] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[14] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[15] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[16] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[17] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[18] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[19] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[1] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[20] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[21] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[22] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[23] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[2] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[3] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[4] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[5] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[6] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[7] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[8] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[9] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.clk ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ena ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[10] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[11] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[12] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[13] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[14] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[15] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[16] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[17] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[1] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[2] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[3] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[4] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[5] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[6] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[7] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[8] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[9] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.k_zero ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[0] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[10] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[11] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[12] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[13] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[14] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[15] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[16] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[17] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[18] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[19] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[1] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[20] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[21] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[22] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[23] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[2] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[3] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[4] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[5] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[6] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[7] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[8] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[9] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.clk ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.ena ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[10] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[11] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[12] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[13] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[14] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[15] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[16] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[17] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[1] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[2] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[3] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[4] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[5] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[6] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[7] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[8] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[9] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.k_zero ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.ow[0] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.ow[10] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.ow[11] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.ow[12] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.ow[13] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.ow[14] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.ow[15] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.ow[16] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.ow[17] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.ow[18] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.ow[19] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.ow[1] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.ow[20] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.ow[21] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.ow[22] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.ow[23] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.ow[2] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.ow[3] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.ow[4] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.ow[5] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.ow[6] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.ow[7] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.ow[8] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.ow[9] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.clk ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ena ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[10] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[11] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[12] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[13] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[14] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[15] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[16] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[17] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[1] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[2] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[3] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[4] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[5] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[6] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[7] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[8] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[9] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.k_zero ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[0] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[10] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[11] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[12] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[13] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[14] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[15] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[16] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[17] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[18] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[19] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[1] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[20] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[21] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[22] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[23] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[2] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[3] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[4] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[5] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[6] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[7] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[8] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[9] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.clk ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ena ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[10] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[11] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[12] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[13] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[14] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[15] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[16] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[17] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[1] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[2] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[3] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[4] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[5] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[6] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[7] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[8] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[9] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.k_zero ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[0] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[10] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[11] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[12] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[13] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[14] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[15] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[16] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[17] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[18] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[19] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[1] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[20] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[21] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[22] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[23] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[2] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[3] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[4] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[5] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[6] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[7] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[8] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[9] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.clk ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ena ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[10] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[11] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[12] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[13] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[14] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[15] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[16] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[17] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[1] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[2] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[3] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[4] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[5] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[6] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[7] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[8] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[9] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.k_zero ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[0] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[10] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[11] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[12] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[13] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[14] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[15] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[16] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[17] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[18] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[19] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[1] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[20] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[21] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[22] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[23] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[2] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[3] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[4] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[5] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[6] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[7] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[8] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[9] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.clk ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.ena ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[10] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[11] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[12] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[13] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[14] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[15] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[16] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[17] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[1] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[2] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[3] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[4] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[5] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[6] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[7] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[8] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[9] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.clk ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ena ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[10] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[11] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[12] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[13] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[14] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[15] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[16] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[17] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[1] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[2] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[3] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[4] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[5] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[6] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[7] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[8] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[9] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.k_zero ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[0] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[10] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[11] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[12] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[13] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[14] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[15] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[16] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[17] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[18] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[19] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[1] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[20] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[21] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[22] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[23] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[2] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[3] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[4] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[5] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[6] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[7] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[8] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[9] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.clk ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.ena ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[10] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[11] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[12] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[13] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[14] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[15] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[16] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[17] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[1] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[2] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[3] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[4] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[5] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[6] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[7] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[8] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[9] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.clk ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ena ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[10] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[11] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[12] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[13] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[14] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[15] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[16] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[17] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[1] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[2] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[3] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[4] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[5] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[6] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[7] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[8] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[9] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.k_zero ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[0] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[10] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[11] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[12] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[13] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[14] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[15] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[16] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[17] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[18] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[19] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[1] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[20] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[21] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[22] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[23] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[2] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[3] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[4] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[5] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[6] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[7] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[8] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[9] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.clk ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.ena ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[10] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[11] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[12] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[13] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[14] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[15] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[16] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[17] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[1] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[2] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[3] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[4] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[5] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[6] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[7] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[8] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[9] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.clk ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ena ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[10] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[11] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[12] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[13] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[14] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[15] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[16] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[17] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[1] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[2] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[3] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[4] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[5] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[6] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[7] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[8] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[9] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.k_zero ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[0] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[10] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[11] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[12] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[13] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[14] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[15] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[16] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[17] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[18] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[19] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[1] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[20] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[21] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[22] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[23] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[2] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[3] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[4] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[5] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[6] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[7] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[8] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[9] ;
 wire \tt_top1.branch[0].l_addr[0] ;
 wire \tt_top1.branch[0].l_k_one ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.clk ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ena ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[10] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[11] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[12] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[13] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[14] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[15] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[16] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[17] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[1] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[2] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[3] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[4] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[5] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[6] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[7] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[8] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[9] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.k_zero ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[0] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[10] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[11] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[12] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[13] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[14] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[15] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[16] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[17] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[18] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[19] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[1] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[20] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[21] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[22] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[23] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[2] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[3] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[4] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[5] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[6] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[7] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[8] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[9] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.clk ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ena ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[10] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[11] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[12] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[13] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[14] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[15] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[16] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[17] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[1] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[2] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[3] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[4] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[5] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[6] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[7] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[8] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[9] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.k_zero ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[0] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[10] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[11] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[12] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[13] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[14] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[15] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[16] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[17] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[18] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[19] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[1] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[20] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[21] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[22] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[23] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[2] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[3] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[4] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[5] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[6] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[7] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[8] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[9] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.clk ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ena ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[10] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[11] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[12] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[13] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[14] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[15] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[16] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[17] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[1] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[2] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[3] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[4] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[5] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[6] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[7] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[8] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[9] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.k_zero ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[0] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[10] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[11] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[12] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[13] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[14] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[15] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[16] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[17] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[18] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[19] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[1] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[20] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[21] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[22] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[23] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[2] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[3] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[4] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[5] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[6] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[7] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[8] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[9] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.clk ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ena ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[10] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[11] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[12] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[13] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[14] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[15] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[16] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[17] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[1] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[2] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[3] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[4] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[5] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[6] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[7] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[8] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[9] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.k_zero ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[0] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[10] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[11] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[12] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[13] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[14] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[15] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[16] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[17] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[18] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[19] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[1] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[20] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[21] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[22] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[23] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[2] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[3] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[4] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[5] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[6] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[7] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[8] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[9] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.clk ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ena ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[10] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[11] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[12] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[13] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[14] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[15] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[16] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[17] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[1] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[2] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[3] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[4] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[5] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[6] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[7] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[8] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[9] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.k_zero ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[0] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[10] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[11] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[12] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[13] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[14] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[15] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[16] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[17] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[18] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[19] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[1] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[20] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[21] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[22] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[23] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[2] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[3] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[4] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[5] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[6] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[7] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[8] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[9] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.clk ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ena ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[10] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[11] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[12] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[13] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[14] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[15] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[16] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[17] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[1] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[2] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[3] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[4] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[5] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[6] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[7] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[8] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[9] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.k_zero ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[0] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[10] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[11] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[12] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[13] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[14] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[15] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[16] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[17] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[18] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[19] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[1] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[20] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[21] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[22] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[23] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[2] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[3] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[4] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[5] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[6] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[7] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[8] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[9] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.clk ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ena ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[10] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[11] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[12] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[13] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[14] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[15] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[16] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[17] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[1] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[2] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[3] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[4] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[5] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[6] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[7] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[8] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[9] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.k_zero ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[0] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[10] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[11] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[12] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[13] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[14] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[15] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[16] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[17] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[18] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[19] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[1] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[20] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[21] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[22] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[23] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[2] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[3] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[4] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[5] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[6] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[7] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[8] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[9] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.clk ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ena ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[10] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[11] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[12] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[13] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[14] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[15] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[16] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[17] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[1] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[2] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[3] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[4] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[5] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[6] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[7] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[8] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[9] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.k_zero ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[0] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[10] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[11] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[12] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[13] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[14] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[15] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[16] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[17] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[18] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[19] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[1] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[20] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[21] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[22] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[23] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[2] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[3] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[4] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[5] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[6] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[7] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[8] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[9] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.clk ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ena ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[10] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[11] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[12] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[13] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[14] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[15] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[16] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[17] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[1] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[2] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[3] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[4] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[5] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[6] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[7] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[8] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[9] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.k_zero ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[0] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[10] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[11] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[12] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[13] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[14] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[15] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[16] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[17] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[18] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[19] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[1] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[20] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[21] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[22] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[23] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[2] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[3] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[4] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[5] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[6] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[7] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[8] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[9] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.clk ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ena ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[10] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[11] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[12] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[13] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[14] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[15] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[16] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[17] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[1] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[2] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[3] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[4] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[5] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[6] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[7] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[8] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[9] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.k_zero ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[0] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[10] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[11] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[12] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[13] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[14] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[15] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[16] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[17] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[18] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[19] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[1] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[20] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[21] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[22] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[23] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[2] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[3] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[4] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[5] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[6] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[7] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[8] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[9] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.clk ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ena ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[10] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[11] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[12] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[13] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[14] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[15] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[16] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[17] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[1] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[2] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[3] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[4] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[5] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[6] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[7] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[8] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[9] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.k_zero ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[0] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[10] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[11] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[12] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[13] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[14] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[15] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[16] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[17] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[18] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[19] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[1] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[20] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[21] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[22] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[23] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[2] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[3] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[4] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[5] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[6] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[7] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[8] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[9] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.clk ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ena ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[10] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[11] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[12] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[13] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[14] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[15] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[16] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[17] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[1] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[2] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[3] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[4] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[5] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[6] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[7] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[8] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[9] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.k_zero ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[0] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[10] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[11] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[12] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[13] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[14] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[15] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[16] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[17] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[18] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[19] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[1] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[20] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[21] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[22] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[23] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[2] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[3] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[4] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[5] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[6] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[7] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[8] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[9] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.clk ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ena ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[10] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[11] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[12] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[13] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[14] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[15] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[16] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[17] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[1] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[2] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[3] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[4] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[5] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[6] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[7] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[8] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[9] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.k_zero ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[0] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[10] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[11] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[12] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[13] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[14] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[15] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[16] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[17] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[18] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[19] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[1] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[20] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[21] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[22] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[23] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[2] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[3] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[4] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[5] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[6] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[7] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[8] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[9] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.clk ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ena ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[10] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[11] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[12] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[13] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[14] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[15] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[16] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[17] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[1] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[2] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[3] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[4] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[5] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[6] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[7] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[8] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[9] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.k_zero ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[0] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[10] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[11] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[12] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[13] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[14] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[15] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[16] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[17] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[18] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[19] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[1] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[20] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[21] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[22] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[23] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[2] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[3] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[4] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[5] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[6] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[7] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[8] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[9] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.clk ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ena ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[10] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[11] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[12] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[13] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[14] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[15] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[16] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[17] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[1] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[2] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[3] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[4] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[5] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[6] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[7] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[8] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[9] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.k_zero ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[0] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[10] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[11] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[12] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[13] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[14] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[15] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[16] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[17] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[18] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[19] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[1] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[20] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[21] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[22] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[23] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[2] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[3] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[4] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[5] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[6] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[7] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[8] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[9] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_addr0[0] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_addr0[1] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_addr0[2] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_addr0[3] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_addr0[4] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_addr0[5] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_addr0[6] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_addr0[7] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_addr0[8] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_clk0 ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_csb0 ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[0] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[10] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[11] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[12] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[13] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[14] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[15] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[16] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[17] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[18] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[19] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[1] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[20] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[21] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[22] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[23] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[24] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[25] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[26] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[27] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[28] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[29] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[2] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[30] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[31] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[3] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[4] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[5] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[6] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[7] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[8] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[9] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[0] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[10] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[11] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[12] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[13] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[14] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[15] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[16] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[17] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[18] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[19] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[1] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[20] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[21] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[22] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[23] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[24] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[25] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[26] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[27] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[28] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[29] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[2] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[30] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[31] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[3] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[4] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[5] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[6] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[7] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[8] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[9] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_web0 ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_wmask0[0] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_wmask0[1] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_wmask0[2] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_wmask0[3] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.clk ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ena ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[10] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[11] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[12] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[13] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[14] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[15] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[16] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[17] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[1] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[2] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[3] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[4] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[5] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[6] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[7] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[8] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[9] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.k_zero ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[0] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[10] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[11] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[12] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[13] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[14] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[15] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[16] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[17] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[18] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[19] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[1] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[20] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[21] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[22] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[23] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[2] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[3] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[4] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[5] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[6] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[7] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[8] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[9] ;
 wire \tt_top1.branch[1].l_addr[0] ;
 wire \tt_top1.branch[1].l_addr[1] ;
 wire \tt_top1.spine_iw[0] ;
 wire \tt_top1.spine_iw[12] ;
 wire \tt_top1.spine_iw[13] ;
 wire \tt_top1.spine_iw[14] ;
 wire \tt_top1.spine_iw[15] ;
 wire \tt_top1.spine_iw[16] ;
 wire \tt_top1.spine_iw[17] ;
 wire \tt_top1.spine_iw[18] ;
 wire \tt_top1.spine_iw[19] ;
 wire \tt_top1.spine_iw[1] ;
 wire \tt_top1.spine_iw[20] ;
 wire \tt_top1.spine_iw[21] ;
 wire \tt_top1.spine_iw[22] ;
 wire \tt_top1.spine_iw[23] ;
 wire \tt_top1.spine_iw[24] ;
 wire \tt_top1.spine_iw[25] ;
 wire \tt_top1.spine_iw[26] ;
 wire \tt_top1.spine_iw[27] ;
 wire \tt_top1.spine_iw[28] ;
 wire \tt_top1.spine_iw[29] ;
 wire \tt_top1.spine_iw[30] ;
 wire \tt_top1.spine_ow[0] ;
 wire \tt_top1.spine_ow[10] ;
 wire \tt_top1.spine_ow[11] ;
 wire \tt_top1.spine_ow[12] ;
 wire \tt_top1.spine_ow[13] ;
 wire \tt_top1.spine_ow[14] ;
 wire \tt_top1.spine_ow[15] ;
 wire \tt_top1.spine_ow[16] ;
 wire \tt_top1.spine_ow[17] ;
 wire \tt_top1.spine_ow[18] ;
 wire \tt_top1.spine_ow[19] ;
 wire \tt_top1.spine_ow[1] ;
 wire \tt_top1.spine_ow[20] ;
 wire \tt_top1.spine_ow[21] ;
 wire \tt_top1.spine_ow[22] ;
 wire \tt_top1.spine_ow[23] ;
 wire \tt_top1.spine_ow[24] ;
 wire \tt_top1.spine_ow[25] ;
 wire \tt_top1.spine_ow[2] ;
 wire \tt_top1.spine_ow[3] ;
 wire \tt_top1.spine_ow[4] ;
 wire \tt_top1.spine_ow[5] ;
 wire \tt_top1.spine_ow[6] ;
 wire \tt_top1.spine_ow[7] ;
 wire \tt_top1.spine_ow[8] ;
 wire \tt_top1.spine_ow[9] ;

 tt_um_as1802 \tt_top1.branch[0].col_um[0].um_bot_I.block_0_0.tt_um_I  (.clk(\tt_top1.branch[0].col_um[0].um_bot_I.clk ),
    .ena(\tt_top1.branch[0].col_um[0].um_bot_I.ena ),
    .rst_n(\tt_top1.branch[0].col_um[0].um_bot_I.iw[1] ),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .ui_in({\tt_top1.branch[0].col_um[0].um_bot_I.iw[9] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[8] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[7] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[6] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[5] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[4] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[3] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[2] }),
    .uio_in({\tt_top1.branch[0].col_um[0].um_bot_I.iw[17] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[16] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[15] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[14] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[13] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[12] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[11] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[10] }),
    .uio_oe({\tt_top1.branch[0].col_um[0].um_bot_I.ow[23] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[22] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[21] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[20] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[19] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[18] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[17] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[16] }),
    .uio_out({\tt_top1.branch[0].col_um[0].um_bot_I.ow[15] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[14] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[13] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[12] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[11] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[10] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[9] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[8] }),
    .uo_out({\tt_top1.branch[0].col_um[0].um_bot_I.ow[7] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[6] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[5] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[4] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[3] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[2] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[1] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[0] }));
 tt_um_loopback \tt_top1.branch[0].col_um[0].um_top_I.block_1_0.tt_um_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .clk(\tt_top1.branch[0].col_um[0].um_top_I.clk ),
    .ena(\tt_top1.branch[0].col_um[0].um_top_I.ena ),
    .rst_n(\tt_top1.branch[0].col_um[0].um_top_I.iw[1] ),
    .ui_in({\tt_top1.branch[0].col_um[0].um_top_I.iw[9] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[8] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[7] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[6] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[5] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[4] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[3] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[2] }),
    .uio_in({\tt_top1.branch[0].col_um[0].um_top_I.iw[17] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[16] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[15] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[14] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[13] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[12] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[11] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[10] }),
    .uio_oe({\tt_top1.branch[0].col_um[0].um_top_I.ow[23] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[22] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[21] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[20] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[19] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[18] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[17] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[16] }),
    .uio_out({\tt_top1.branch[0].col_um[0].um_top_I.ow[15] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[14] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[13] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[12] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[11] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[10] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[9] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[8] }),
    .uo_out({\tt_top1.branch[0].col_um[0].um_top_I.ow[7] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[6] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[5] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[4] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[3] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[2] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[1] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[0] }));
 tt_um_urish_simon \tt_top1.branch[0].col_um[1].um_bot_I.block_0_1.tt_um_I  (.clk(\tt_top1.branch[0].col_um[1].um_bot_I.clk ),
    .ena(\tt_top1.branch[0].col_um[1].um_bot_I.ena ),
    .rst_n(\tt_top1.branch[0].col_um[1].um_bot_I.iw[1] ),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .ui_in({\tt_top1.branch[0].col_um[1].um_bot_I.iw[9] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[8] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[7] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[6] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[5] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[4] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[3] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[2] }),
    .uio_in({\tt_top1.branch[0].col_um[1].um_bot_I.iw[17] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[16] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[15] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[14] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[13] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[12] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[11] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[10] }),
    .uio_oe({\tt_top1.branch[0].col_um[1].um_bot_I.ow[23] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[22] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[21] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[20] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[19] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[18] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[17] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[16] }),
    .uio_out({\tt_top1.branch[0].col_um[1].um_bot_I.ow[15] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[14] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[13] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[12] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[11] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[10] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[9] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[8] }),
    .uo_out({\tt_top1.branch[0].col_um[1].um_bot_I.ow[7] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[6] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[5] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[4] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[3] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[2] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[1] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[0] }));
 tt_um_power_test \tt_top1.branch[0].col_um[1].um_top_I.block_1_1.tt_um_I  (.clk(\tt_top1.branch[0].col_um[1].um_top_I.clk ),
    .ena(\tt_top1.branch[0].col_um[1].um_top_I.ena ),
    .rst_n(\tt_top1.branch[0].col_um[1].um_top_I.iw[1] ),
    .vssd1(vssd1),
    .vccd1(vccd1),
    .ui_in({\tt_top1.branch[0].col_um[1].um_top_I.iw[9] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[8] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[7] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[6] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[5] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[4] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[3] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[2] }),
    .uio_in({\tt_top1.branch[0].col_um[1].um_top_I.iw[17] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[16] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[15] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[14] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[13] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[12] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[11] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[10] }),
    .uio_oe({\tt_top1.branch[0].col_um[1].um_top_I.ow[23] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[22] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[21] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[20] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[19] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[18] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[17] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[16] }),
    .uio_out({\tt_top1.branch[0].col_um[1].um_top_I.ow[15] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[14] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[13] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[12] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[11] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[10] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[9] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[8] }),
    .uo_out({\tt_top1.branch[0].col_um[1].um_top_I.ow[7] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[6] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[5] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[4] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[3] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[2] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[1] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[0] }));
 tt_um_kiwih_tt_top \tt_top1.branch[0].col_um[2].um_bot_I.block_0_2.tt_um_I  (.clk(\tt_top1.branch[0].col_um[2].um_bot_I.clk ),
    .ena(\tt_top1.branch[0].col_um[2].um_bot_I.ena ),
    .rst_n(\tt_top1.branch[0].col_um[2].um_bot_I.iw[1] ),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .ui_in({\tt_top1.branch[0].col_um[2].um_bot_I.iw[9] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[8] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[7] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[6] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[5] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[4] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[3] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[2] }),
    .uio_in({\tt_top1.branch[0].col_um[2].um_bot_I.iw[17] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[16] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[15] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[14] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[13] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[12] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[11] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[10] }),
    .uio_oe({\tt_top1.branch[0].col_um[2].um_bot_I.ow[23] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[22] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[21] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[20] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[19] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[18] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[17] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[16] }),
    .uio_out({\tt_top1.branch[0].col_um[2].um_bot_I.ow[15] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[14] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[13] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[12] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[11] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[10] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[9] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[8] }),
    .uo_out({\tt_top1.branch[0].col_um[2].um_bot_I.ow[7] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[6] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[5] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[4] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[3] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[2] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[1] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[0] }));
 tt_um_htfab_totp \tt_top1.branch[0].col_um[2].um_top_I.block_1_2.tt_um_I  (.clk(\tt_top1.branch[0].col_um[2].um_top_I.clk ),
    .ena(\tt_top1.branch[0].col_um[2].um_top_I.ena ),
    .rst_n(\tt_top1.branch[0].col_um[2].um_top_I.iw[1] ),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .ui_in({\tt_top1.branch[0].col_um[2].um_top_I.iw[9] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[8] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[7] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[6] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[5] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[4] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[3] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[2] }),
    .uio_in({\tt_top1.branch[0].col_um[2].um_top_I.iw[17] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[16] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[15] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[14] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[13] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[12] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[11] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[10] }),
    .uio_oe({\tt_top1.branch[0].col_um[2].um_top_I.ow[23] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[22] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[21] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[20] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[19] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[18] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[17] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[16] }),
    .uio_out({\tt_top1.branch[0].col_um[2].um_top_I.ow[15] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[14] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[13] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[12] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[11] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[10] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[9] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[8] }),
    .uo_out({\tt_top1.branch[0].col_um[2].um_top_I.ow[7] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[6] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[5] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[4] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[3] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[2] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[1] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[0] }));
 tt_um_wokwi_366318576852367361 \tt_top1.branch[0].col_um[3].um_bot_I.block_0_3.tt_um_I  (.clk(\tt_top1.branch[0].col_um[3].um_bot_I.clk ),
    .ena(\tt_top1.branch[0].col_um[3].um_bot_I.ena ),
    .rst_n(\tt_top1.branch[0].col_um[3].um_bot_I.iw[1] ),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .ui_in({\tt_top1.branch[0].col_um[3].um_bot_I.iw[9] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[8] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[7] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[6] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[5] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[4] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[3] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[2] }),
    .uio_in({\tt_top1.branch[0].col_um[3].um_bot_I.iw[17] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[16] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[15] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[14] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[13] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[12] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[11] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[10] }),
    .uio_oe({\tt_top1.branch[0].col_um[3].um_bot_I.ow[23] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[22] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[21] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[20] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[19] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[18] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[17] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[16] }),
    .uio_out({\tt_top1.branch[0].col_um[3].um_bot_I.ow[15] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[14] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[13] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[12] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[11] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[10] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[9] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[8] }),
    .uo_out({\tt_top1.branch[0].col_um[3].um_bot_I.ow[7] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[6] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[5] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[4] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[3] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[2] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[1] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[0] }));
 tt_um_gatecat_fpga_top \tt_top1.branch[0].col_um[3].um_top_I.block_1_3.tt_um_I  (.clk(\tt_top1.branch[0].col_um[3].um_top_I.clk ),
    .ena(\tt_top1.branch[0].col_um[3].um_top_I.ena ),
    .rst_n(\tt_top1.branch[0].col_um[3].um_top_I.iw[1] ),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .ui_in({\tt_top1.branch[0].col_um[3].um_top_I.iw[9] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[8] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[7] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[6] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[5] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[4] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[3] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[2] }),
    .uio_in({\tt_top1.branch[0].col_um[3].um_top_I.iw[17] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[16] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[15] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[14] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[13] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[12] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[11] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[10] }),
    .uio_oe({\tt_top1.branch[0].col_um[3].um_top_I.ow[23] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[22] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[21] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[20] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[19] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[18] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[17] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[16] }),
    .uio_out({\tt_top1.branch[0].col_um[3].um_top_I.ow[15] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[14] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[13] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[12] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[11] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[10] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[9] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[8] }),
    .uo_out({\tt_top1.branch[0].col_um[3].um_top_I.ow[7] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[6] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[5] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[4] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[3] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[2] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[1] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[0] }));
 tt_um_urish_dffram \tt_top1.branch[0].col_um[4].um_bot_I.block_0_4.tt_um_I  (.clk(\tt_top1.branch[0].col_um[4].um_bot_I.clk ),
    .ena(\tt_top1.branch[0].col_um[4].um_bot_I.ena ),
    .rst_n(\tt_top1.branch[0].col_um[4].um_bot_I.iw[1] ),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .ui_in({\tt_top1.branch[0].col_um[4].um_bot_I.iw[9] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[8] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[7] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[6] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[5] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[4] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[3] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[2] }),
    .uio_in({\tt_top1.branch[0].col_um[4].um_bot_I.iw[17] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[16] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[15] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[14] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[13] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[12] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[11] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[10] }),
    .uio_oe({\tt_top1.branch[0].col_um[4].um_bot_I.ow[23] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[22] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[21] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[20] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[19] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[18] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[17] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[16] }),
    .uio_out({\tt_top1.branch[0].col_um[4].um_bot_I.ow[15] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[14] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[13] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[12] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[11] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[10] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[9] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[8] }),
    .uo_out({\tt_top1.branch[0].col_um[4].um_bot_I.ow[7] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[6] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[5] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[4] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[3] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[2] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[1] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[0] }));
 tt_um_Reloj_top \tt_top1.branch[0].col_um[4].um_top_I.block_1_4.tt_um_I  (.clk(\tt_top1.branch[0].col_um[4].um_top_I.clk ),
    .ena(\tt_top1.branch[0].col_um[4].um_top_I.ena ),
    .rst_n(\tt_top1.branch[0].col_um[4].um_top_I.iw[1] ),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .ui_in({\tt_top1.branch[0].col_um[4].um_top_I.iw[9] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[8] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[7] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[6] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[5] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[4] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[3] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[2] }),
    .uio_in({\tt_top1.branch[0].col_um[4].um_top_I.iw[17] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[16] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[15] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[14] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[13] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[12] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[11] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[10] }),
    .uio_oe({\tt_top1.branch[0].col_um[4].um_top_I.ow[23] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[22] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[21] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[20] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[19] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[18] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[17] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[16] }),
    .uio_out({\tt_top1.branch[0].col_um[4].um_top_I.ow[15] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[14] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[13] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[12] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[11] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[10] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[9] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[8] }),
    .uo_out({\tt_top1.branch[0].col_um[4].um_top_I.ow[7] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[6] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[5] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[4] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[3] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[2] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[1] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[0] }));
 tt_um_algofoogle_solo_squash \tt_top1.branch[0].col_um[5].um_top_I.block_1_5.tt_um_I  (.clk(\tt_top1.branch[0].col_um[5].um_top_I.clk ),
    .ena(\tt_top1.branch[0].col_um[5].um_top_I.ena ),
    .rst_n(\tt_top1.branch[0].col_um[5].um_top_I.iw[1] ),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .ui_in({\tt_top1.branch[0].col_um[5].um_top_I.iw[9] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[8] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[7] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[6] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[5] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[4] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[3] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[2] }),
    .uio_in({\tt_top1.branch[0].col_um[5].um_top_I.iw[17] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[16] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[15] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[14] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[13] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[12] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[11] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[10] }),
    .uio_oe({\tt_top1.branch[0].col_um[5].um_top_I.ow[23] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[22] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[21] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[20] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[19] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[18] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[17] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[16] }),
    .uio_out({\tt_top1.branch[0].col_um[5].um_top_I.ow[15] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[14] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[13] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[12] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[11] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[10] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[9] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[8] }),
    .uo_out({\tt_top1.branch[0].col_um[5].um_top_I.ow[7] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[6] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[5] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[4] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[3] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[2] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[1] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[0] }));
 tt_um_apu_pulse \tt_top1.branch[0].col_um[6].um_top_I.block_1_6.tt_um_I  (.clk(\tt_top1.branch[0].col_um[6].um_top_I.clk ),
    .ena(\tt_top1.branch[0].col_um[6].um_top_I.ena ),
    .rst_n(\tt_top1.branch[0].col_um[6].um_top_I.iw[1] ),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .ui_in({\tt_top1.branch[0].col_um[6].um_top_I.iw[9] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[8] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[7] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[6] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[5] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[4] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[3] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[2] }),
    .uio_in({\tt_top1.branch[0].col_um[6].um_top_I.iw[17] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[16] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[15] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[14] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[13] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[12] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[11] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[10] }),
    .uio_oe({\tt_top1.branch[0].col_um[6].um_top_I.ow[23] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[22] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[21] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[20] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[19] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[18] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[17] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[16] }),
    .uio_out({\tt_top1.branch[0].col_um[6].um_top_I.ow[15] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[14] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[13] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[12] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[11] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[10] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[9] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[8] }),
    .uo_out({\tt_top1.branch[0].col_um[6].um_top_I.ow[7] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[6] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[5] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[4] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[3] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[2] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[1] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[0] }));
 tt_um_thorkn_vgaclock \tt_top1.branch[0].col_um[7].um_top_I.block_1_7.tt_um_I  (.clk(\tt_top1.branch[0].col_um[7].um_top_I.clk ),
    .ena(\tt_top1.branch[0].col_um[7].um_top_I.ena ),
    .rst_n(\tt_top1.branch[0].col_um[7].um_top_I.iw[1] ),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .ui_in({\tt_top1.branch[0].col_um[7].um_top_I.iw[9] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[8] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[7] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[6] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[5] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[4] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[3] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[2] }),
    .uio_in({\tt_top1.branch[0].col_um[7].um_top_I.iw[17] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[16] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[15] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[14] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[13] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[12] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[11] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[10] }),
    .uio_oe({\tt_top1.branch[0].col_um[7].um_top_I.ow[23] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[22] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[21] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[20] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[19] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[18] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[17] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[16] }),
    .uio_out({\tt_top1.branch[0].col_um[7].um_top_I.ow[15] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[14] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[13] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[12] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[11] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[10] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[9] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[8] }),
    .uo_out({\tt_top1.branch[0].col_um[7].um_top_I.ow[7] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[6] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[5] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[4] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[3] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[2] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[1] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[0] }));
 tt_mux \tt_top1.branch[0].mux_I  (.k_one(\tt_top1.branch[0].l_k_one ),
    .k_zero(\tt_top1.branch[0].l_addr[0] ),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .addr({\tt_top1.branch[0].l_addr[0] ,
    \tt_top1.branch[0].l_addr[0] ,
    \tt_top1.branch[0].l_addr[0] ,
    \tt_top1.branch[0].l_addr[0] ,
    \tt_top1.branch[0].l_addr[0] }),
    .spine_iw({\tt_top1.spine_iw[30] ,
    \tt_top1.spine_iw[29] ,
    \tt_top1.spine_iw[28] ,
    \tt_top1.spine_iw[27] ,
    \tt_top1.spine_iw[26] ,
    \tt_top1.spine_iw[25] ,
    \tt_top1.spine_iw[24] ,
    \tt_top1.spine_iw[23] ,
    \tt_top1.spine_iw[22] ,
    \tt_top1.spine_iw[21] ,
    \tt_top1.spine_iw[20] ,
    \tt_top1.spine_iw[19] ,
    \tt_top1.spine_iw[18] ,
    \tt_top1.spine_iw[17] ,
    \tt_top1.spine_iw[16] ,
    \tt_top1.spine_iw[15] ,
    \tt_top1.spine_iw[14] ,
    \tt_top1.spine_iw[13] ,
    \tt_top1.spine_iw[12] ,
    la_data_out[9],
    la_data_out[8],
    la_data_out[7],
    la_data_out[6],
    la_data_out[5],
    la_data_out[4],
    la_data_out[3],
    la_data_out[2],
    la_data_out[1],
    la_data_out[0],
    \tt_top1.spine_iw[1] ,
    \tt_top1.spine_iw[0] }),
    .spine_ow({\tt_top1.spine_ow[25] ,
    \tt_top1.spine_ow[24] ,
    \tt_top1.spine_ow[23] ,
    \tt_top1.spine_ow[22] ,
    \tt_top1.spine_ow[21] ,
    \tt_top1.spine_ow[20] ,
    \tt_top1.spine_ow[19] ,
    \tt_top1.spine_ow[18] ,
    \tt_top1.spine_ow[17] ,
    \tt_top1.spine_ow[16] ,
    \tt_top1.spine_ow[15] ,
    \tt_top1.spine_ow[14] ,
    \tt_top1.spine_ow[13] ,
    \tt_top1.spine_ow[12] ,
    \tt_top1.spine_ow[11] ,
    \tt_top1.spine_ow[10] ,
    \tt_top1.spine_ow[9] ,
    \tt_top1.spine_ow[8] ,
    \tt_top1.spine_ow[7] ,
    \tt_top1.spine_ow[6] ,
    \tt_top1.spine_ow[5] ,
    \tt_top1.spine_ow[4] ,
    \tt_top1.spine_ow[3] ,
    \tt_top1.spine_ow[2] ,
    \tt_top1.spine_ow[1] ,
    \tt_top1.spine_ow[0] }),
    .um_ena({\tt_top1.branch[0].col_um[7].um_top_I.ena ,
    \tt_top1.branch[0].col_um[7].um_bot_I.ena ,
    \tt_top1.branch[0].col_um[6].um_top_I.ena ,
    \tt_top1.branch[0].col_um[6].um_bot_I.ena ,
    \tt_top1.branch[0].col_um[5].um_top_I.ena ,
    \tt_top1.branch[0].col_um[5].um_bot_I.ena ,
    \tt_top1.branch[0].col_um[4].um_top_I.ena ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ena ,
    \tt_top1.branch[0].col_um[3].um_top_I.ena ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ena ,
    \tt_top1.branch[0].col_um[2].um_top_I.ena ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ena ,
    \tt_top1.branch[0].col_um[1].um_top_I.ena ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ena ,
    \tt_top1.branch[0].col_um[0].um_top_I.ena ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ena }),
    .um_iw({\tt_top1.branch[0].col_um[7].um_top_I.iw[17] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[16] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[15] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[14] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[13] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[12] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[11] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[10] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[9] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[8] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[7] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[6] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[5] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[4] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[3] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[2] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[1] ,
    \tt_top1.branch[0].col_um[7].um_top_I.clk ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[17] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[16] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[15] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[14] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[13] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[12] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[11] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[10] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[9] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[8] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[7] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[6] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[5] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[4] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[3] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[2] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[1] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.clk ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[17] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[16] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[15] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[14] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[13] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[12] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[11] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[10] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[9] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[8] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[7] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[6] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[5] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[4] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[3] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[2] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[1] ,
    \tt_top1.branch[0].col_um[6].um_top_I.clk ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[17] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[16] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[15] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[14] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[13] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[12] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[11] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[10] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[9] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[8] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[7] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[6] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[5] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[4] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[3] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[2] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[1] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.clk ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[17] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[16] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[15] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[14] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[13] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[12] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[11] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[10] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[9] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[8] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[7] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[6] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[5] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[4] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[3] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[2] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[1] ,
    \tt_top1.branch[0].col_um[5].um_top_I.clk ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[17] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[16] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[15] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[14] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[13] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[12] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[11] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[10] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[9] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[8] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[7] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[6] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[5] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[4] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[3] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[2] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[1] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.clk ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[17] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[16] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[15] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[14] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[13] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[12] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[11] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[10] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[9] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[8] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[7] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[6] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[5] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[4] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[3] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[2] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[1] ,
    \tt_top1.branch[0].col_um[4].um_top_I.clk ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[17] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[16] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[15] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[14] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[13] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[12] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[11] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[10] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[9] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[8] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[7] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[6] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[5] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[4] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[3] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[2] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[1] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.clk ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[17] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[16] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[15] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[14] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[13] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[12] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[11] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[10] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[9] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[8] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[7] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[6] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[5] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[4] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[3] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[2] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[1] ,
    \tt_top1.branch[0].col_um[3].um_top_I.clk ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[17] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[16] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[15] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[14] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[13] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[12] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[11] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[10] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[9] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[8] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[7] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[6] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[5] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[4] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[3] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[2] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[1] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.clk ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[17] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[16] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[15] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[14] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[13] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[12] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[11] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[10] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[9] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[8] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[7] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[6] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[5] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[4] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[3] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[2] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[1] ,
    \tt_top1.branch[0].col_um[2].um_top_I.clk ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[17] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[16] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[15] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[14] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[13] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[12] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[11] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[10] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[9] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[8] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[7] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[6] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[5] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[4] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[3] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[2] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[1] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.clk ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[17] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[16] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[15] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[14] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[13] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[12] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[11] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[10] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[9] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[8] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[7] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[6] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[5] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[4] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[3] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[2] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[1] ,
    \tt_top1.branch[0].col_um[1].um_top_I.clk ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[17] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[16] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[15] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[14] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[13] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[12] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[11] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[10] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[9] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[8] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[7] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[6] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[5] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[4] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[3] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[2] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[1] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.clk ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[17] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[16] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[15] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[14] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[13] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[12] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[11] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[10] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[9] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[8] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[7] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[6] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[5] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[4] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[3] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[2] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[1] ,
    \tt_top1.branch[0].col_um[0].um_top_I.clk ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[17] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[16] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[15] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[14] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[13] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[12] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[11] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[10] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[9] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[8] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[7] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[6] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[5] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[4] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[3] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[2] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[1] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.clk }),
    .um_k_zero({\tt_top1.branch[0].col_um[7].um_top_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_top_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_top_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[4].um_top_I.k_zero ,
    \tt_top1.branch[0].col_um[4].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[3].um_top_I.k_zero ,
    \tt_top1.branch[0].col_um[3].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[2].um_top_I.k_zero ,
    \tt_top1.branch[0].col_um[2].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[1].um_top_I.k_zero ,
    \tt_top1.branch[0].col_um[1].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[0].um_top_I.k_zero ,
    \tt_top1.branch[0].col_um[0].um_bot_I.k_zero }),
    .um_ow({\tt_top1.branch[0].col_um[7].um_top_I.ow[23] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[22] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[21] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[20] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[19] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[18] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[17] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[16] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[15] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[14] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[13] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[12] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[11] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[10] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[9] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[8] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[7] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[6] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[5] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[4] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[3] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[2] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[1] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[0] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[23] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[22] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[21] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[20] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[19] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[18] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[17] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[16] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[15] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[14] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[13] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[12] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[11] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[10] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[9] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[8] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[7] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[6] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[5] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[4] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[3] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[2] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[1] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[0] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[23] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[22] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[21] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[20] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[19] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[18] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[17] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[16] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[15] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[14] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[13] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[12] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[11] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[10] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[9] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[8] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[7] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[6] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[5] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[4] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[3] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[2] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[1] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[0] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[23] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[22] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[21] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[20] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[19] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[18] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[17] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[16] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[15] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[14] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[13] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[12] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[11] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[10] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[9] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[8] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[7] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[6] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[5] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[4] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[3] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[2] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[1] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[0] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[23] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[22] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[21] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[20] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[19] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[18] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[17] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[16] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[15] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[14] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[13] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[12] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[11] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[10] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[9] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[8] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[7] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[6] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[5] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[4] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[3] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[2] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[1] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[0] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[23] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[22] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[21] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[20] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[19] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[18] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[17] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[16] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[15] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[14] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[13] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[12] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[11] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[10] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[9] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[8] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[7] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[6] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[5] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[4] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[3] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[2] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[1] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[0] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[23] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[22] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[21] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[20] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[19] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[18] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[17] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[16] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[15] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[14] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[13] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[12] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[11] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[10] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[9] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[8] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[7] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[6] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[5] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[4] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[3] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[2] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[1] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ow[0] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[23] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[22] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[21] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[20] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[19] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[18] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[17] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[16] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[15] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[14] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[13] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[12] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[11] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[10] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[9] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[8] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[7] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[6] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[5] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[4] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[3] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[2] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[1] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[0] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[23] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[22] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[21] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[20] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[19] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[18] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[17] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[16] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[15] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[14] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[13] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[12] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[11] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[10] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[9] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[8] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[7] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[6] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[5] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[4] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[3] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[2] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[1] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[0] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[23] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[22] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[21] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[20] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[19] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[18] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[17] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[16] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[15] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[14] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[13] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[12] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[11] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[10] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[9] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[8] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[7] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[6] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[5] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[4] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[3] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[2] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[1] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[0] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[23] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[22] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[21] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[20] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[19] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[18] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[17] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[16] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[15] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[14] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[13] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[12] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[11] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[10] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[9] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[8] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[7] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[6] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[5] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[4] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[3] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[2] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[1] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[0] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[23] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[22] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[21] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[20] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[19] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[18] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[17] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[16] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[15] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[14] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[13] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[12] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[11] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[10] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[9] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[8] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[7] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[6] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[5] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[4] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[3] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[2] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[1] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[0] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[23] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[22] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[21] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[20] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[19] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[18] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[17] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[16] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[15] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[14] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[13] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[12] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[11] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[10] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[9] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[8] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[7] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[6] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[5] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[4] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[3] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[2] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[1] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[0] }));
 tt_um_greycode_top \tt_top1.branch[1].col_um[0].um_bot_I.block_0_16.tt_um_I  (.clk(\tt_top1.branch[1].col_um[0].um_bot_I.clk ),
    .ena(\tt_top1.branch[1].col_um[0].um_bot_I.ena ),
    .rst_n(\tt_top1.branch[1].col_um[0].um_bot_I.iw[1] ),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .ui_in({\tt_top1.branch[1].col_um[0].um_bot_I.iw[9] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[8] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[7] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[6] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[5] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[4] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[3] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[2] }),
    .uio_in({\tt_top1.branch[1].col_um[0].um_bot_I.iw[17] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[16] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[15] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[14] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[13] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[12] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[11] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[10] }),
    .uio_oe({\tt_top1.branch[1].col_um[0].um_bot_I.ow[23] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[22] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[21] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[20] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[19] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[18] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[17] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[16] }),
    .uio_out({\tt_top1.branch[1].col_um[0].um_bot_I.ow[15] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[14] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[13] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[12] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[11] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[10] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[9] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[8] }),
    .uo_out({\tt_top1.branch[1].col_um[0].um_bot_I.ow[7] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[6] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[5] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[4] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[3] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[2] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[1] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[0] }));
 tt_um_ringosc_cnt_pfet \tt_top1.branch[1].col_um[0].um_top_I.block_1_16.tt_um_I  (.clk(\tt_top1.branch[1].col_um[0].um_top_I.clk ),
    .ena(\tt_top1.branch[1].col_um[0].um_top_I.ena ),
    .rst_n(\tt_top1.branch[1].col_um[0].um_top_I.iw[1] ),
    .vssd1(vssd1),
    .vccd1(vccd1),
    .ui_in({\tt_top1.branch[1].col_um[0].um_top_I.iw[9] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[8] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[7] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[6] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[5] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[4] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[3] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[2] }),
    .uio_in({\tt_top1.branch[1].col_um[0].um_top_I.iw[17] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[16] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[15] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[14] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[13] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[12] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[11] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[10] }),
    .uio_oe({\tt_top1.branch[1].col_um[0].um_top_I.ow[23] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[22] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[21] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[20] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[19] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[18] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[17] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[16] }),
    .uio_out({\tt_top1.branch[1].col_um[0].um_top_I.ow[15] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[14] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[13] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[12] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[11] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[10] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[9] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[8] }),
    .uo_out({\tt_top1.branch[1].col_um[0].um_top_I.ow[7] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[6] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[5] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[4] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[3] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[2] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[1] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[0] }));
 tt_um_moyes0_top_module \tt_top1.branch[1].col_um[1].um_bot_I.block_0_17.tt_um_I  (.clk(\tt_top1.branch[1].col_um[1].um_bot_I.clk ),
    .ena(\tt_top1.branch[1].col_um[1].um_bot_I.ena ),
    .rst_n(\tt_top1.branch[1].col_um[1].um_bot_I.iw[1] ),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .ui_in({\tt_top1.branch[1].col_um[1].um_bot_I.iw[9] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[8] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[7] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[6] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[5] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[4] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[3] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[2] }),
    .uio_in({\tt_top1.branch[1].col_um[1].um_bot_I.iw[17] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[16] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[15] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[14] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[13] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[12] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[11] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[10] }),
    .uio_oe({\tt_top1.branch[1].col_um[1].um_bot_I.ow[23] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[22] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[21] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[20] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[19] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[18] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[17] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[16] }),
    .uio_out({\tt_top1.branch[1].col_um[1].um_bot_I.ow[15] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[14] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[13] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[12] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[11] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[10] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[9] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[8] }),
    .uo_out({\tt_top1.branch[1].col_um[1].um_bot_I.ow[7] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[6] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[5] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[4] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[3] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[2] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[1] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[0] }));
 tt_um_wokwi_347497504164545108 \tt_top1.branch[1].col_um[1].um_top_I.block_1_17.tt_um_I  (.clk(\tt_top1.branch[1].col_um[1].um_top_I.clk ),
    .ena(\tt_top1.branch[1].col_um[1].um_top_I.ena ),
    .rst_n(\tt_top1.branch[1].col_um[1].um_top_I.iw[1] ),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .ui_in({\tt_top1.branch[1].col_um[1].um_top_I.iw[9] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[8] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[7] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[6] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[5] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[4] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[3] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[2] }),
    .uio_in({\tt_top1.branch[1].col_um[1].um_top_I.iw[17] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[16] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[15] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[14] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[13] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[12] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[11] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[10] }),
    .uio_oe({\tt_top1.branch[1].col_um[1].um_top_I.ow[23] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[22] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[21] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[20] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[19] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[18] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[17] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[16] }),
    .uio_out({\tt_top1.branch[1].col_um[1].um_top_I.ow[15] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[14] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[13] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[12] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[11] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[10] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[9] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[8] }),
    .uo_out({\tt_top1.branch[1].col_um[1].um_top_I.ow[7] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[6] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[5] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[4] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[3] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[2] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[1] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[0] }));
 tt_um_vga_clock \tt_top1.branch[1].col_um[2].um_bot_I.block_0_18.tt_um_I  (.clk(\tt_top1.branch[1].col_um[2].um_bot_I.clk ),
    .ena(\tt_top1.branch[1].col_um[2].um_bot_I.ena ),
    .rst_n(\tt_top1.branch[1].col_um[2].um_bot_I.iw[1] ),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .ui_in({\tt_top1.branch[1].col_um[2].um_bot_I.iw[9] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[8] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[7] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[6] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[5] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[4] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[3] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[2] }),
    .uio_in({\tt_top1.branch[1].col_um[2].um_bot_I.iw[17] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[16] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[15] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[14] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[13] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[12] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[11] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[10] }),
    .uio_oe({\tt_top1.branch[1].col_um[2].um_bot_I.ow[23] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[22] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[21] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[20] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[19] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[18] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[17] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[16] }),
    .uio_out({\tt_top1.branch[1].col_um[2].um_bot_I.ow[15] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[14] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[13] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[12] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[11] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[10] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[9] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[8] }),
    .uo_out({\tt_top1.branch[1].col_um[2].um_bot_I.ow[7] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[6] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[5] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[4] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[3] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[2] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[1] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[0] }));
 tt_um_wokwi_347144898258928211 \tt_top1.branch[1].col_um[2].um_top_I.block_1_18.tt_um_I  (.clk(\tt_top1.branch[1].col_um[2].um_top_I.clk ),
    .ena(\tt_top1.branch[1].col_um[2].um_top_I.ena ),
    .rst_n(\tt_top1.branch[1].col_um[2].um_top_I.iw[1] ),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .ui_in({\tt_top1.branch[1].col_um[2].um_top_I.iw[9] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[8] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[7] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[6] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[5] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[4] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[3] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[2] }),
    .uio_in({\tt_top1.branch[1].col_um[2].um_top_I.iw[17] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[16] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[15] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[14] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[13] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[12] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[11] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[10] }),
    .uio_oe({\tt_top1.branch[1].col_um[2].um_top_I.ow[23] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[22] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[21] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[20] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[19] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[18] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[17] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[16] }),
    .uio_out({\tt_top1.branch[1].col_um[2].um_top_I.ow[15] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[14] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[13] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[12] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[11] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[10] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[9] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[8] }),
    .uo_out({\tt_top1.branch[1].col_um[2].um_top_I.ow[7] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[6] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[5] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[4] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[3] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[2] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[1] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[0] }));
 tt_um_TrainLED2_top \tt_top1.branch[1].col_um[3].um_bot_I.block_0_19.tt_um_I  (.clk(\tt_top1.branch[1].col_um[3].um_bot_I.clk ),
    .ena(\tt_top1.branch[1].col_um[3].um_bot_I.ena ),
    .rst_n(\tt_top1.branch[1].col_um[3].um_bot_I.iw[1] ),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .ui_in({\tt_top1.branch[1].col_um[3].um_bot_I.iw[9] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[8] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[7] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[6] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[5] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[4] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[3] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[2] }),
    .uio_in({\tt_top1.branch[1].col_um[3].um_bot_I.iw[17] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[16] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[15] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[14] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[13] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[12] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[11] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[10] }),
    .uio_oe({\tt_top1.branch[1].col_um[3].um_bot_I.ow[23] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[22] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[21] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[20] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[19] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[18] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[17] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[16] }),
    .uio_out({\tt_top1.branch[1].col_um[3].um_bot_I.ow[15] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[14] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[13] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[12] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[11] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[10] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[9] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[8] }),
    .uo_out({\tt_top1.branch[1].col_um[3].um_bot_I.ow[7] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[6] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[5] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[4] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[3] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[2] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[1] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[0] }));
 tt_um_wokwi_347417602591556180 \tt_top1.branch[1].col_um[3].um_top_I.block_1_19.tt_um_I  (.clk(\tt_top1.branch[1].col_um[3].um_top_I.clk ),
    .ena(\tt_top1.branch[1].col_um[3].um_top_I.ena ),
    .rst_n(\tt_top1.branch[1].col_um[3].um_top_I.iw[1] ),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .ui_in({\tt_top1.branch[1].col_um[3].um_top_I.iw[9] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[8] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[7] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[6] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[5] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[4] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[3] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[2] }),
    .uio_in({\tt_top1.branch[1].col_um[3].um_top_I.iw[17] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[16] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[15] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[14] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[13] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[12] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[11] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[10] }),
    .uio_oe({\tt_top1.branch[1].col_um[3].um_top_I.ow[23] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[22] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[21] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[20] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[19] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[18] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[17] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[16] }),
    .uio_out({\tt_top1.branch[1].col_um[3].um_top_I.ow[15] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[14] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[13] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[12] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[11] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[10] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[9] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[8] }),
    .uo_out({\tt_top1.branch[1].col_um[3].um_top_I.ow[7] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[6] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[5] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[4] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[3] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[2] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[1] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[0] }));
 tt_um_tomkeddie_a \tt_top1.branch[1].col_um[4].um_bot_I.block_0_20.tt_um_I  (.clk(\tt_top1.branch[1].col_um[4].um_bot_I.clk ),
    .ena(\tt_top1.branch[1].col_um[4].um_bot_I.ena ),
    .rst_n(\tt_top1.branch[1].col_um[4].um_bot_I.iw[1] ),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .ui_in({\tt_top1.branch[1].col_um[4].um_bot_I.iw[9] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[8] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[7] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[6] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[5] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[4] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[3] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[2] }),
    .uio_in({\tt_top1.branch[1].col_um[4].um_bot_I.iw[17] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[16] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[15] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[14] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[13] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[12] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[11] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[10] }),
    .uio_oe({\tt_top1.branch[1].col_um[4].um_bot_I.ow[23] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[22] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[21] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[20] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[19] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[18] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[17] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[16] }),
    .uio_out({\tt_top1.branch[1].col_um[4].um_bot_I.ow[15] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[14] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[13] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[12] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[11] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[10] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[9] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[8] }),
    .uo_out({\tt_top1.branch[1].col_um[4].um_bot_I.ow[7] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[6] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[5] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[4] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[3] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[2] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[1] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[0] }));
 tt_um_millerresearch_top \tt_top1.branch[1].col_um[4].um_top_I.block_1_20.tt_um_I  (.clk(\tt_top1.branch[1].col_um[4].um_top_I.clk ),
    .ena(\tt_top1.branch[1].col_um[4].um_top_I.ena ),
    .rst_n(\tt_top1.branch[1].col_um[4].um_top_I.iw[1] ),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .ui_in({\tt_top1.branch[1].col_um[4].um_top_I.iw[9] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[8] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[7] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[6] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[5] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[4] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[3] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[2] }),
    .uio_in({\tt_top1.branch[1].col_um[4].um_top_I.iw[17] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[16] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[15] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[14] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[13] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[12] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[11] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[10] }),
    .uio_oe({\tt_top1.branch[1].col_um[4].um_top_I.ow[23] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[22] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[21] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[20] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[19] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[18] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[17] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[16] }),
    .uio_out({\tt_top1.branch[1].col_um[4].um_top_I.ow[15] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[14] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[13] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[12] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[11] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[10] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[9] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[8] }),
    .uo_out({\tt_top1.branch[1].col_um[4].um_top_I.ow[7] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[6] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[5] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[4] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[3] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[2] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[1] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[0] }));
 tt_um_ternaryPC_radixconvert \tt_top1.branch[1].col_um[5].um_bot_I.block_0_21.tt_um_I  (.clk(\tt_top1.branch[1].col_um[5].um_bot_I.clk ),
    .ena(\tt_top1.branch[1].col_um[5].um_bot_I.ena ),
    .rst_n(\tt_top1.branch[1].col_um[5].um_bot_I.iw[1] ),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .ui_in({\tt_top1.branch[1].col_um[5].um_bot_I.iw[9] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[8] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[7] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[6] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[5] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[4] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[3] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[2] }),
    .uio_in({\tt_top1.branch[1].col_um[5].um_bot_I.iw[17] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[16] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[15] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[14] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[13] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[12] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[11] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[10] }),
    .uio_oe({\tt_top1.branch[1].col_um[5].um_bot_I.ow[23] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[22] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[21] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[20] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[19] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[18] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[17] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[16] }),
    .uio_out({\tt_top1.branch[1].col_um[5].um_bot_I.ow[15] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[14] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[13] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[12] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[11] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[10] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[9] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[8] }),
    .uo_out({\tt_top1.branch[1].col_um[5].um_bot_I.ow[7] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[6] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[5] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[4] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[3] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[2] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[1] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[0] }));
 tt_um_psychogenic_neptuneproportional \tt_top1.branch[1].col_um[5].um_top_I.block_1_21.tt_um_I  (.clk(\tt_top1.branch[1].col_um[5].um_top_I.clk ),
    .ena(\tt_top1.branch[1].col_um[5].um_top_I.ena ),
    .rst_n(\tt_top1.branch[1].col_um[5].um_top_I.iw[1] ),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .ui_in({\tt_top1.branch[1].col_um[5].um_top_I.iw[9] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[8] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[7] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[6] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[5] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[4] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[3] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[2] }),
    .uio_in({\tt_top1.branch[1].col_um[5].um_top_I.iw[17] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[16] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[15] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[14] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[13] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[12] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[11] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[10] }),
    .uio_oe({\tt_top1.branch[1].col_um[5].um_top_I.ow[23] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[22] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[21] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[20] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[19] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[18] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[17] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[16] }),
    .uio_out({\tt_top1.branch[1].col_um[5].um_top_I.ow[15] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[14] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[13] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[12] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[11] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[10] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[9] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[8] }),
    .uo_out({\tt_top1.branch[1].col_um[5].um_top_I.ow[7] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[6] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[5] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[4] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[3] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[2] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[1] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[0] }));
 tt_um_MichaelBell_hovalaag \tt_top1.branch[1].col_um[6].um_bot_I.block_0_22.tt_um_I  (.clk(\tt_top1.branch[1].col_um[6].um_bot_I.clk ),
    .ena(\tt_top1.branch[1].col_um[6].um_bot_I.ena ),
    .rst_n(\tt_top1.branch[1].col_um[6].um_bot_I.iw[1] ),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .ui_in({\tt_top1.branch[1].col_um[6].um_bot_I.iw[9] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[8] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[7] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[6] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[5] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[4] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[3] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[2] }),
    .uio_in({\tt_top1.branch[1].col_um[6].um_bot_I.iw[17] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[16] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[15] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[14] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[13] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[12] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[11] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[10] }),
    .uio_oe({\tt_top1.branch[1].col_um[6].um_bot_I.ow[23] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[22] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[21] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[20] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[19] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[18] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[17] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[16] }),
    .uio_out({\tt_top1.branch[1].col_um[6].um_bot_I.ow[15] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[14] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[13] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[12] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[11] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[10] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[9] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[8] }),
    .uo_out({\tt_top1.branch[1].col_um[6].um_bot_I.ow[7] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[6] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[5] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[4] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[3] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[2] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[1] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[0] }));
 tt_um_test \tt_top1.branch[1].col_um[6].um_top_I.block_1_22.tt_um_I  (.clk(\tt_top1.branch[1].col_um[6].um_top_I.clk ),
    .ena(\tt_top1.branch[1].col_um[6].um_top_I.ena ),
    .rst_n(\tt_top1.branch[1].col_um[6].um_top_I.iw[1] ),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .ui_in({\tt_top1.branch[1].col_um[6].um_top_I.iw[9] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[8] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[7] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[6] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[5] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[4] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[3] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[2] }),
    .uio_in({\tt_top1.branch[1].col_um[6].um_top_I.iw[17] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[16] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[15] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[14] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[13] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[12] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[11] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[10] }),
    .uio_oe({\tt_top1.branch[1].col_um[6].um_top_I.ow[23] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[22] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[21] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[20] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[19] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[18] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[17] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[16] }),
    .uio_out({\tt_top1.branch[1].col_um[6].um_top_I.ow[15] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[14] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[13] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[12] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[11] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[10] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[9] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[8] }),
    .uo_out({\tt_top1.branch[1].col_um[6].um_top_I.ow[7] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[6] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[5] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[4] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[3] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[2] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[1] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[0] }));
 tt_um_cam \tt_top1.branch[1].col_um[7].um_bot_I.block_0_23.tt_um_I  (.clk(\tt_top1.branch[1].col_um[7].um_bot_I.clk ),
    .ena(\tt_top1.branch[1].col_um[7].um_bot_I.ena ),
    .rst_n(\tt_top1.branch[1].col_um[7].um_bot_I.iw[1] ),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .ui_in({\tt_top1.branch[1].col_um[7].um_bot_I.iw[9] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[8] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[7] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[6] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[5] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[4] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[3] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[2] }),
    .uio_in({\tt_top1.branch[1].col_um[7].um_bot_I.iw[17] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[16] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[15] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[14] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[13] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[12] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[11] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[10] }),
    .uio_oe({\tt_top1.branch[1].col_um[7].um_bot_I.ow[23] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[22] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[21] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[20] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[19] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[18] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[17] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[16] }),
    .uio_out({\tt_top1.branch[1].col_um[7].um_bot_I.ow[15] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[14] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[13] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[12] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[11] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[10] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[9] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[8] }),
    .uo_out({\tt_top1.branch[1].col_um[7].um_bot_I.ow[7] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[6] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[5] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[4] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[3] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[2] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[1] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[0] }));
 sky130_sram_2kbyte_1rw1r_32x512_8 \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.sram  (.csb0(\tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_csb0 ),
    .csb1(\tt_top1.branch[1].col_um[7].um_top_I.k_zero ),
    .web0(\tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_web0 ),
    .clk0(\tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_clk0 ),
    .clk1(\tt_top1.branch[1].col_um[7].um_top_I.k_zero ),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .addr0({\tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_addr0[8] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_addr0[7] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_addr0[6] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_addr0[5] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_addr0[4] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_addr0[3] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_addr0[2] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_addr0[1] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_addr0[0] }),
    .addr1({\tt_top1.branch[1].col_um[7].um_top_I.k_zero ,
    \tt_top1.branch[1].col_um[7].um_top_I.k_zero ,
    \tt_top1.branch[1].col_um[7].um_top_I.k_zero ,
    \tt_top1.branch[1].col_um[7].um_top_I.k_zero ,
    \tt_top1.branch[1].col_um[7].um_top_I.k_zero ,
    \tt_top1.branch[1].col_um[7].um_top_I.k_zero ,
    \tt_top1.branch[1].col_um[7].um_top_I.k_zero ,
    \tt_top1.branch[1].col_um[7].um_top_I.k_zero ,
    \tt_top1.branch[1].col_um[7].um_top_I.k_zero }),
    .din0({\tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[31] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[30] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[29] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[28] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[27] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[26] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[25] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[24] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[23] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[22] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[21] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[20] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[19] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[18] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[17] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[16] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[15] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[14] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[13] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[12] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[11] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[10] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[9] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[8] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[7] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[6] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[5] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[4] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[3] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[2] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[1] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[0] }),
    .dout0({\tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[31] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[30] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[29] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[28] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[27] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[26] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[25] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[24] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[23] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[22] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[21] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[20] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[19] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[18] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[17] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[16] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[15] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[14] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[13] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[12] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[11] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[10] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[9] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[8] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[7] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[6] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[5] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[4] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[3] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[2] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[1] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[0] }),
    .dout1({_NC1,
    _NC2,
    _NC3,
    _NC4,
    _NC5,
    _NC6,
    _NC7,
    _NC8,
    _NC9,
    _NC10,
    _NC11,
    _NC12,
    _NC13,
    _NC14,
    _NC15,
    _NC16,
    _NC17,
    _NC18,
    _NC19,
    _NC20,
    _NC21,
    _NC22,
    _NC23,
    _NC24,
    _NC25,
    _NC26,
    _NC27,
    _NC28,
    _NC29,
    _NC30,
    _NC31,
    _NC32}),
    .wmask0({\tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_wmask0[3] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_wmask0[2] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_wmask0[1] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_wmask0[0] }));
 tt_um_urish_sram_poc \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.tt_um_I  (.clk(\tt_top1.branch[1].col_um[7].um_top_I.clk ),
    .ena(\tt_top1.branch[1].col_um[7].um_top_I.ena ),
    .ram_clk0(\tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_clk0 ),
    .ram_csb0(\tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_csb0 ),
    .ram_web0(\tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_web0 ),
    .rst_n(\tt_top1.branch[1].col_um[7].um_top_I.iw[1] ),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .ram_addr0({\tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_addr0[8] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_addr0[7] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_addr0[6] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_addr0[5] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_addr0[4] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_addr0[3] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_addr0[2] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_addr0[1] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_addr0[0] }),
    .ram_din0({\tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[31] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[30] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[29] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[28] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[27] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[26] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[25] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[24] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[23] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[22] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[21] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[20] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[19] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[18] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[17] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[16] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[15] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[14] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[13] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[12] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[11] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[10] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[9] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[8] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[7] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[6] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[5] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[4] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[3] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[2] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[1] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_din0[0] }),
    .ram_dout0({\tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[31] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[30] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[29] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[28] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[27] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[26] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[25] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[24] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[23] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[22] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[21] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[20] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[19] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[18] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[17] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[16] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[15] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[14] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[13] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[12] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[11] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[10] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[9] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[8] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[7] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[6] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[5] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[4] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[3] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[2] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[1] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_dout0[0] }),
    .ram_wmask0({\tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_wmask0[3] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_wmask0[2] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_wmask0[1] ,
    \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.ram_wmask0[0] }),
    .ui_in({\tt_top1.branch[1].col_um[7].um_top_I.iw[9] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[8] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[7] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[6] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[5] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[4] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[3] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[2] }),
    .uio_in({\tt_top1.branch[1].col_um[7].um_top_I.iw[17] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[16] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[15] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[14] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[13] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[12] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[11] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[10] }),
    .uio_oe({\tt_top1.branch[1].col_um[7].um_top_I.ow[23] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[22] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[21] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[20] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[19] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[18] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[17] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[16] }),
    .uio_out({\tt_top1.branch[1].col_um[7].um_top_I.ow[15] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[14] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[13] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[12] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[11] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[10] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[9] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[8] }),
    .uo_out({\tt_top1.branch[1].col_um[7].um_top_I.ow[7] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[6] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[5] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[4] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[3] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[2] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[1] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[0] }));
 tt_mux \tt_top1.branch[1].mux_I  (.k_one(\tt_top1.branch[1].l_addr[0] ),
    .k_zero(\tt_top1.branch[1].l_addr[1] ),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .addr({\tt_top1.branch[1].l_addr[1] ,
    \tt_top1.branch[1].l_addr[1] ,
    \tt_top1.branch[1].l_addr[1] ,
    \tt_top1.branch[1].l_addr[1] ,
    \tt_top1.branch[1].l_addr[0] }),
    .spine_iw({\tt_top1.spine_iw[30] ,
    \tt_top1.spine_iw[29] ,
    \tt_top1.spine_iw[28] ,
    \tt_top1.spine_iw[27] ,
    \tt_top1.spine_iw[26] ,
    \tt_top1.spine_iw[25] ,
    \tt_top1.spine_iw[24] ,
    \tt_top1.spine_iw[23] ,
    \tt_top1.spine_iw[22] ,
    \tt_top1.spine_iw[21] ,
    \tt_top1.spine_iw[20] ,
    \tt_top1.spine_iw[19] ,
    \tt_top1.spine_iw[18] ,
    \tt_top1.spine_iw[17] ,
    \tt_top1.spine_iw[16] ,
    \tt_top1.spine_iw[15] ,
    \tt_top1.spine_iw[14] ,
    \tt_top1.spine_iw[13] ,
    \tt_top1.spine_iw[12] ,
    la_data_out[9],
    la_data_out[8],
    la_data_out[7],
    la_data_out[6],
    la_data_out[5],
    la_data_out[4],
    la_data_out[3],
    la_data_out[2],
    la_data_out[1],
    la_data_out[0],
    \tt_top1.spine_iw[1] ,
    \tt_top1.spine_iw[0] }),
    .spine_ow({\tt_top1.spine_ow[25] ,
    \tt_top1.spine_ow[24] ,
    \tt_top1.spine_ow[23] ,
    \tt_top1.spine_ow[22] ,
    \tt_top1.spine_ow[21] ,
    \tt_top1.spine_ow[20] ,
    \tt_top1.spine_ow[19] ,
    \tt_top1.spine_ow[18] ,
    \tt_top1.spine_ow[17] ,
    \tt_top1.spine_ow[16] ,
    \tt_top1.spine_ow[15] ,
    \tt_top1.spine_ow[14] ,
    \tt_top1.spine_ow[13] ,
    \tt_top1.spine_ow[12] ,
    \tt_top1.spine_ow[11] ,
    \tt_top1.spine_ow[10] ,
    \tt_top1.spine_ow[9] ,
    \tt_top1.spine_ow[8] ,
    \tt_top1.spine_ow[7] ,
    \tt_top1.spine_ow[6] ,
    \tt_top1.spine_ow[5] ,
    \tt_top1.spine_ow[4] ,
    \tt_top1.spine_ow[3] ,
    \tt_top1.spine_ow[2] ,
    \tt_top1.spine_ow[1] ,
    \tt_top1.spine_ow[0] }),
    .um_ena({\tt_top1.branch[1].col_um[7].um_top_I.ena ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ena ,
    \tt_top1.branch[1].col_um[6].um_top_I.ena ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ena ,
    \tt_top1.branch[1].col_um[5].um_top_I.ena ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ena ,
    \tt_top1.branch[1].col_um[4].um_top_I.ena ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ena ,
    \tt_top1.branch[1].col_um[3].um_top_I.ena ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ena ,
    \tt_top1.branch[1].col_um[2].um_top_I.ena ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ena ,
    \tt_top1.branch[1].col_um[1].um_top_I.ena ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ena ,
    \tt_top1.branch[1].col_um[0].um_top_I.ena ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ena }),
    .um_iw({\tt_top1.branch[1].col_um[7].um_top_I.iw[17] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[16] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[15] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[14] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[13] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[12] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[11] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[10] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[9] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[8] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[7] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[6] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[5] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[4] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[3] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[2] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[1] ,
    \tt_top1.branch[1].col_um[7].um_top_I.clk ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[17] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[16] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[15] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[14] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[13] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[12] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[11] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[10] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[9] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[8] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[7] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[6] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[5] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[4] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[3] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[2] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[1] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.clk ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[17] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[16] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[15] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[14] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[13] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[12] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[11] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[10] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[9] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[8] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[7] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[6] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[5] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[4] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[3] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[2] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[1] ,
    \tt_top1.branch[1].col_um[6].um_top_I.clk ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[17] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[16] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[15] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[14] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[13] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[12] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[11] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[10] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[9] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[8] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[7] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[6] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[5] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[4] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[3] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[2] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[1] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.clk ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[17] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[16] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[15] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[14] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[13] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[12] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[11] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[10] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[9] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[8] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[7] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[6] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[5] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[4] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[3] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[2] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[1] ,
    \tt_top1.branch[1].col_um[5].um_top_I.clk ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[17] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[16] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[15] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[14] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[13] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[12] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[11] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[10] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[9] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[8] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[7] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[6] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[5] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[4] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[3] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[2] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[1] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.clk ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[17] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[16] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[15] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[14] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[13] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[12] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[11] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[10] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[9] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[8] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[7] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[6] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[5] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[4] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[3] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[2] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[1] ,
    \tt_top1.branch[1].col_um[4].um_top_I.clk ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[17] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[16] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[15] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[14] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[13] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[12] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[11] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[10] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[9] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[8] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[7] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[6] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[5] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[4] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[3] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[2] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[1] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.clk ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[17] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[16] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[15] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[14] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[13] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[12] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[11] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[10] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[9] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[8] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[7] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[6] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[5] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[4] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[3] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[2] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[1] ,
    \tt_top1.branch[1].col_um[3].um_top_I.clk ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[17] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[16] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[15] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[14] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[13] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[12] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[11] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[10] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[9] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[8] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[7] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[6] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[5] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[4] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[3] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[2] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[1] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.clk ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[17] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[16] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[15] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[14] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[13] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[12] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[11] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[10] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[9] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[8] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[7] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[6] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[5] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[4] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[3] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[2] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[1] ,
    \tt_top1.branch[1].col_um[2].um_top_I.clk ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[17] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[16] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[15] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[14] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[13] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[12] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[11] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[10] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[9] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[8] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[7] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[6] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[5] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[4] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[3] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[2] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[1] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.clk ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[17] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[16] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[15] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[14] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[13] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[12] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[11] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[10] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[9] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[8] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[7] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[6] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[5] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[4] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[3] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[2] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[1] ,
    \tt_top1.branch[1].col_um[1].um_top_I.clk ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[17] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[16] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[15] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[14] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[13] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[12] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[11] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[10] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[9] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[8] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[7] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[6] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[5] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[4] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[3] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[2] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[1] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.clk ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[17] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[16] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[15] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[14] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[13] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[12] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[11] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[10] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[9] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[8] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[7] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[6] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[5] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[4] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[3] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[2] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[1] ,
    \tt_top1.branch[1].col_um[0].um_top_I.clk ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[17] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[16] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[15] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[14] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[13] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[12] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[11] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[10] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[9] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[8] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[7] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[6] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[5] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[4] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[3] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[2] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[1] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.clk }),
    .um_k_zero({\tt_top1.branch[1].col_um[7].um_top_I.k_zero ,
    \tt_top1.branch[1].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[1].col_um[6].um_top_I.k_zero ,
    \tt_top1.branch[1].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[1].col_um[5].um_top_I.k_zero ,
    \tt_top1.branch[1].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[1].col_um[4].um_top_I.k_zero ,
    \tt_top1.branch[1].col_um[4].um_bot_I.k_zero ,
    \tt_top1.branch[1].col_um[3].um_top_I.k_zero ,
    \tt_top1.branch[1].col_um[3].um_bot_I.k_zero ,
    \tt_top1.branch[1].col_um[2].um_top_I.k_zero ,
    \tt_top1.branch[1].col_um[2].um_bot_I.k_zero ,
    \tt_top1.branch[1].col_um[1].um_top_I.k_zero ,
    \tt_top1.branch[1].col_um[1].um_bot_I.k_zero ,
    \tt_top1.branch[1].col_um[0].um_top_I.k_zero ,
    \tt_top1.branch[1].col_um[0].um_bot_I.k_zero }),
    .um_ow({\tt_top1.branch[1].col_um[7].um_top_I.ow[23] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[22] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[21] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[20] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[19] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[18] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[17] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[16] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[15] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[14] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[13] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[12] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[11] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[10] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[9] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[8] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[7] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[6] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[5] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[4] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[3] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[2] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[1] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[0] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[23] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[22] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[21] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[20] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[19] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[18] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[17] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[16] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[15] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[14] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[13] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[12] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[11] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[10] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[9] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[8] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[7] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[6] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[5] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[4] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[3] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[2] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[1] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[0] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[23] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[22] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[21] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[20] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[19] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[18] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[17] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[16] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[15] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[14] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[13] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[12] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[11] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[10] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[9] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[8] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[7] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[6] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[5] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[4] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[3] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[2] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[1] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[0] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[23] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[22] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[21] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[20] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[19] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[18] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[17] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[16] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[15] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[14] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[13] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[12] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[11] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[10] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[9] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[8] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[7] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[6] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[5] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[4] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[3] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[2] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[1] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[0] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[23] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[22] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[21] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[20] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[19] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[18] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[17] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[16] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[15] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[14] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[13] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[12] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[11] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[10] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[9] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[8] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[7] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[6] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[5] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[4] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[3] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[2] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[1] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[0] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[23] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[22] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[21] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[20] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[19] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[18] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[17] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[16] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[15] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[14] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[13] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[12] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[11] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[10] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[9] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[8] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[7] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[6] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[5] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[4] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[3] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[2] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[1] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[0] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[23] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[22] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[21] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[20] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[19] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[18] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[17] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[16] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[15] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[14] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[13] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[12] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[11] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[10] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[9] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[8] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[7] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[6] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[5] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[4] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[3] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[2] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[1] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[0] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[23] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[22] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[21] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[20] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[19] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[18] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[17] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[16] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[15] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[14] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[13] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[12] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[11] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[10] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[9] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[8] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[7] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[6] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[5] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[4] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[3] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[2] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[1] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[0] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[23] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[22] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[21] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[20] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[19] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[18] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[17] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[16] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[15] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[14] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[13] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[12] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[11] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[10] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[9] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[8] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[7] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[6] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[5] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[4] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[3] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[2] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[1] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[0] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[23] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[22] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[21] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[20] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[19] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[18] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[17] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[16] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[15] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[14] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[13] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[12] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[11] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[10] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[9] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[8] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[7] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[6] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[5] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[4] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[3] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[2] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[1] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[0] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[23] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[22] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[21] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[20] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[19] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[18] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[17] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[16] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[15] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[14] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[13] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[12] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[11] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[10] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[9] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[8] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[7] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[6] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[5] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[4] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[3] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[2] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[1] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[0] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[23] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[22] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[21] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[20] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[19] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[18] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[17] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[16] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[15] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[14] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[13] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[12] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[11] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[10] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[9] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[8] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[7] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[6] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[5] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[4] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[3] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[2] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[1] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[0] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[23] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[22] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[21] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[20] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[19] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[18] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[17] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[16] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[15] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[14] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[13] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[12] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[11] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[10] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[9] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[8] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[7] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[6] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[5] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[4] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[3] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[2] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[1] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[0] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[23] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[22] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[21] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[20] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[19] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[18] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[17] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[16] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[15] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[14] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[13] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[12] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[11] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[10] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[9] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[8] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[7] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[6] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[5] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[4] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[3] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[2] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[1] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[0] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[23] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[22] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[21] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[20] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[19] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[18] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[17] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[16] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[15] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[14] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[13] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[12] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[11] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[10] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[9] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[8] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[7] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[6] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[5] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[4] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[3] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[2] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[1] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[0] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[23] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[22] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[21] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[20] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[19] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[18] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[17] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[16] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[15] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[14] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[13] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[12] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[11] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[10] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[9] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[8] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[7] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[6] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[5] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[4] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[3] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[2] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[1] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[0] }));
 tt_ctrl \tt_top1.ctrl_I  (.ctrl_ena(io_in[32]),
    .ctrl_sel_inc(io_in[34]),
    .ctrl_sel_rst_n(io_in[36]),
    .k_one(\tt_top1.io_oeb[0] ),
    .k_zero(wbs_ack_o),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .pad_ui_in({io_in[15],
    io_in[14],
    io_in[13],
    io_in[12],
    io_in[11],
    io_in[10],
    io_in[9],
    io_in[8],
    io_in[7],
    io_in[6]}),
    .pad_uio_in({io_in[31],
    io_in[30],
    io_in[29],
    io_in[28],
    io_in[27],
    io_in[26],
    io_in[25],
    io_in[24]}),
    .pad_uio_oe_n({io_oeb[31],
    io_oeb[30],
    io_oeb[29],
    io_oeb[28],
    io_oeb[27],
    io_oeb[26],
    io_oeb[25],
    io_oeb[24]}),
    .pad_uio_out({io_out[31],
    io_out[30],
    io_out[29],
    io_out[28],
    io_out[27],
    io_out[26],
    io_out[25],
    io_out[24]}),
    .pad_uo_out({io_out[23],
    io_out[22],
    io_out[21],
    io_out[20],
    io_out[19],
    io_out[18],
    io_out[17],
    io_out[16]}),
    .spine_iw({\tt_top1.spine_iw[30] ,
    \tt_top1.spine_iw[29] ,
    \tt_top1.spine_iw[28] ,
    \tt_top1.spine_iw[27] ,
    \tt_top1.spine_iw[26] ,
    \tt_top1.spine_iw[25] ,
    \tt_top1.spine_iw[24] ,
    \tt_top1.spine_iw[23] ,
    \tt_top1.spine_iw[22] ,
    \tt_top1.spine_iw[21] ,
    \tt_top1.spine_iw[20] ,
    \tt_top1.spine_iw[19] ,
    \tt_top1.spine_iw[18] ,
    \tt_top1.spine_iw[17] ,
    \tt_top1.spine_iw[16] ,
    \tt_top1.spine_iw[15] ,
    \tt_top1.spine_iw[14] ,
    \tt_top1.spine_iw[13] ,
    \tt_top1.spine_iw[12] ,
    la_data_out[9],
    la_data_out[8],
    la_data_out[7],
    la_data_out[6],
    la_data_out[5],
    la_data_out[4],
    la_data_out[3],
    la_data_out[2],
    la_data_out[1],
    la_data_out[0],
    \tt_top1.spine_iw[1] ,
    \tt_top1.spine_iw[0] }),
    .spine_ow({\tt_top1.spine_ow[25] ,
    \tt_top1.spine_ow[24] ,
    \tt_top1.spine_ow[23] ,
    \tt_top1.spine_ow[22] ,
    \tt_top1.spine_ow[21] ,
    \tt_top1.spine_ow[20] ,
    \tt_top1.spine_ow[19] ,
    \tt_top1.spine_ow[18] ,
    \tt_top1.spine_ow[17] ,
    \tt_top1.spine_ow[16] ,
    \tt_top1.spine_ow[15] ,
    \tt_top1.spine_ow[14] ,
    \tt_top1.spine_ow[13] ,
    \tt_top1.spine_ow[12] ,
    \tt_top1.spine_ow[11] ,
    \tt_top1.spine_ow[10] ,
    \tt_top1.spine_ow[9] ,
    \tt_top1.spine_ow[8] ,
    \tt_top1.spine_ow[7] ,
    \tt_top1.spine_ow[6] ,
    \tt_top1.spine_ow[5] ,
    \tt_top1.spine_ow[4] ,
    \tt_top1.spine_ow[3] ,
    \tt_top1.spine_ow[2] ,
    \tt_top1.spine_ow[1] ,
    \tt_top1.spine_ow[0] }));
 assign io_oeb[0] = \tt_top1.io_oeb[0] ;
 assign io_oeb[10] = \tt_top1.io_oeb[0] ;
 assign io_oeb[11] = \tt_top1.io_oeb[0] ;
 assign io_oeb[12] = \tt_top1.io_oeb[0] ;
 assign io_oeb[13] = \tt_top1.io_oeb[0] ;
 assign io_oeb[14] = \tt_top1.io_oeb[0] ;
 assign io_oeb[15] = \tt_top1.io_oeb[0] ;
 assign io_oeb[16] = wbs_ack_o;
 assign io_oeb[17] = wbs_ack_o;
 assign io_oeb[18] = wbs_ack_o;
 assign io_oeb[19] = wbs_ack_o;
 assign io_oeb[1] = \tt_top1.io_oeb[0] ;
 assign io_oeb[20] = wbs_ack_o;
 assign io_oeb[21] = wbs_ack_o;
 assign io_oeb[22] = wbs_ack_o;
 assign io_oeb[23] = wbs_ack_o;
 assign io_oeb[2] = \tt_top1.io_oeb[0] ;
 assign io_oeb[32] = \tt_top1.io_oeb[0] ;
 assign io_oeb[33] = wbs_ack_o;
 assign io_oeb[34] = \tt_top1.io_oeb[0] ;
 assign io_oeb[35] = wbs_ack_o;
 assign io_oeb[36] = \tt_top1.io_oeb[0] ;
 assign io_oeb[37] = wbs_ack_o;
 assign io_oeb[3] = \tt_top1.io_oeb[0] ;
 assign io_oeb[4] = wbs_ack_o;
 assign io_oeb[5] = wbs_ack_o;
 assign io_oeb[6] = \tt_top1.io_oeb[0] ;
 assign io_oeb[7] = \tt_top1.io_oeb[0] ;
 assign io_oeb[8] = \tt_top1.io_oeb[0] ;
 assign io_oeb[9] = \tt_top1.io_oeb[0] ;
 assign io_out[0] = \tt_top1.io_oeb[0] ;
 assign io_out[10] = \tt_top1.io_oeb[0] ;
 assign io_out[11] = \tt_top1.io_oeb[0] ;
 assign io_out[12] = \tt_top1.io_oeb[0] ;
 assign io_out[13] = \tt_top1.io_oeb[0] ;
 assign io_out[14] = \tt_top1.io_oeb[0] ;
 assign io_out[15] = \tt_top1.io_oeb[0] ;
 assign io_out[1] = \tt_top1.io_oeb[0] ;
 assign io_out[2] = \tt_top1.io_oeb[0] ;
 assign io_out[32] = wbs_ack_o;
 assign io_out[33] = wbs_ack_o;
 assign io_out[34] = wbs_ack_o;
 assign io_out[35] = wbs_ack_o;
 assign io_out[36] = wbs_ack_o;
 assign io_out[37] = wbs_ack_o;
 assign io_out[3] = \tt_top1.io_oeb[0] ;
 assign io_out[4] = wbs_ack_o;
 assign io_out[5] = user_clock2;
 assign io_out[6] = \tt_top1.io_oeb[0] ;
 assign io_out[7] = \tt_top1.io_oeb[0] ;
 assign io_out[8] = \tt_top1.io_oeb[0] ;
 assign io_out[9] = \tt_top1.io_oeb[0] ;
 assign la_data_out[100] = wbs_ack_o;
 assign la_data_out[101] = wbs_ack_o;
 assign la_data_out[102] = wbs_ack_o;
 assign la_data_out[103] = wbs_ack_o;
 assign la_data_out[104] = wbs_ack_o;
 assign la_data_out[105] = wbs_ack_o;
 assign la_data_out[106] = wbs_ack_o;
 assign la_data_out[107] = wbs_ack_o;
 assign la_data_out[108] = wbs_ack_o;
 assign la_data_out[109] = wbs_ack_o;
 assign la_data_out[10] = wbs_ack_o;
 assign la_data_out[110] = wbs_ack_o;
 assign la_data_out[111] = wbs_ack_o;
 assign la_data_out[112] = wbs_ack_o;
 assign la_data_out[113] = wbs_ack_o;
 assign la_data_out[114] = wbs_ack_o;
 assign la_data_out[115] = wbs_ack_o;
 assign la_data_out[116] = wbs_ack_o;
 assign la_data_out[117] = wbs_ack_o;
 assign la_data_out[118] = wbs_ack_o;
 assign la_data_out[119] = wbs_ack_o;
 assign la_data_out[11] = wbs_ack_o;
 assign la_data_out[120] = wbs_ack_o;
 assign la_data_out[121] = wbs_ack_o;
 assign la_data_out[122] = wbs_ack_o;
 assign la_data_out[123] = wbs_ack_o;
 assign la_data_out[124] = wbs_ack_o;
 assign la_data_out[125] = wbs_ack_o;
 assign la_data_out[126] = wbs_ack_o;
 assign la_data_out[127] = wbs_ack_o;
 assign la_data_out[12] = wbs_ack_o;
 assign la_data_out[13] = wbs_ack_o;
 assign la_data_out[14] = wbs_ack_o;
 assign la_data_out[15] = wbs_ack_o;
 assign la_data_out[16] = wbs_ack_o;
 assign la_data_out[17] = wbs_ack_o;
 assign la_data_out[18] = wbs_ack_o;
 assign la_data_out[19] = wbs_ack_o;
 assign la_data_out[20] = wbs_ack_o;
 assign la_data_out[21] = wbs_ack_o;
 assign la_data_out[22] = wbs_ack_o;
 assign la_data_out[23] = wbs_ack_o;
 assign la_data_out[24] = wbs_ack_o;
 assign la_data_out[25] = wbs_ack_o;
 assign la_data_out[26] = wbs_ack_o;
 assign la_data_out[27] = wbs_ack_o;
 assign la_data_out[28] = wbs_ack_o;
 assign la_data_out[29] = wbs_ack_o;
 assign la_data_out[30] = wbs_ack_o;
 assign la_data_out[31] = wbs_ack_o;
 assign la_data_out[32] = wbs_ack_o;
 assign la_data_out[33] = wbs_ack_o;
 assign la_data_out[34] = wbs_ack_o;
 assign la_data_out[35] = wbs_ack_o;
 assign la_data_out[36] = wbs_ack_o;
 assign la_data_out[37] = wbs_ack_o;
 assign la_data_out[38] = wbs_ack_o;
 assign la_data_out[39] = wbs_ack_o;
 assign la_data_out[40] = wbs_ack_o;
 assign la_data_out[41] = wbs_ack_o;
 assign la_data_out[42] = wbs_ack_o;
 assign la_data_out[43] = wbs_ack_o;
 assign la_data_out[44] = wbs_ack_o;
 assign la_data_out[45] = wbs_ack_o;
 assign la_data_out[46] = wbs_ack_o;
 assign la_data_out[47] = wbs_ack_o;
 assign la_data_out[48] = wbs_ack_o;
 assign la_data_out[49] = wbs_ack_o;
 assign la_data_out[50] = wbs_ack_o;
 assign la_data_out[51] = wbs_ack_o;
 assign la_data_out[52] = wbs_ack_o;
 assign la_data_out[53] = wbs_ack_o;
 assign la_data_out[54] = wbs_ack_o;
 assign la_data_out[55] = wbs_ack_o;
 assign la_data_out[56] = wbs_ack_o;
 assign la_data_out[57] = wbs_ack_o;
 assign la_data_out[58] = wbs_ack_o;
 assign la_data_out[59] = wbs_ack_o;
 assign la_data_out[60] = wbs_ack_o;
 assign la_data_out[61] = wbs_ack_o;
 assign la_data_out[62] = wbs_ack_o;
 assign la_data_out[63] = wbs_ack_o;
 assign la_data_out[64] = wbs_ack_o;
 assign la_data_out[65] = wbs_ack_o;
 assign la_data_out[66] = wbs_ack_o;
 assign la_data_out[67] = wbs_ack_o;
 assign la_data_out[68] = wbs_ack_o;
 assign la_data_out[69] = wbs_ack_o;
 assign la_data_out[70] = wbs_ack_o;
 assign la_data_out[71] = wbs_ack_o;
 assign la_data_out[72] = wbs_ack_o;
 assign la_data_out[73] = wbs_ack_o;
 assign la_data_out[74] = wbs_ack_o;
 assign la_data_out[75] = wbs_ack_o;
 assign la_data_out[76] = wbs_ack_o;
 assign la_data_out[77] = wbs_ack_o;
 assign la_data_out[78] = wbs_ack_o;
 assign la_data_out[79] = wbs_ack_o;
 assign la_data_out[80] = wbs_ack_o;
 assign la_data_out[81] = wbs_ack_o;
 assign la_data_out[82] = wbs_ack_o;
 assign la_data_out[83] = wbs_ack_o;
 assign la_data_out[84] = wbs_ack_o;
 assign la_data_out[85] = wbs_ack_o;
 assign la_data_out[86] = wbs_ack_o;
 assign la_data_out[87] = wbs_ack_o;
 assign la_data_out[88] = wbs_ack_o;
 assign la_data_out[89] = wbs_ack_o;
 assign la_data_out[90] = wbs_ack_o;
 assign la_data_out[91] = wbs_ack_o;
 assign la_data_out[92] = wbs_ack_o;
 assign la_data_out[93] = wbs_ack_o;
 assign la_data_out[94] = wbs_ack_o;
 assign la_data_out[95] = wbs_ack_o;
 assign la_data_out[96] = wbs_ack_o;
 assign la_data_out[97] = wbs_ack_o;
 assign la_data_out[98] = wbs_ack_o;
 assign la_data_out[99] = wbs_ack_o;
 assign user_irq[0] = wbs_ack_o;
 assign user_irq[1] = wbs_ack_o;
 assign user_irq[2] = wbs_ack_o;
 assign wbs_dat_o[0] = wbs_ack_o;
 assign wbs_dat_o[10] = wbs_ack_o;
 assign wbs_dat_o[11] = wbs_ack_o;
 assign wbs_dat_o[12] = wbs_ack_o;
 assign wbs_dat_o[13] = wbs_ack_o;
 assign wbs_dat_o[14] = wbs_ack_o;
 assign wbs_dat_o[15] = wbs_ack_o;
 assign wbs_dat_o[16] = wbs_ack_o;
 assign wbs_dat_o[17] = wbs_ack_o;
 assign wbs_dat_o[18] = wbs_ack_o;
 assign wbs_dat_o[19] = wbs_ack_o;
 assign wbs_dat_o[1] = wbs_ack_o;
 assign wbs_dat_o[20] = wbs_ack_o;
 assign wbs_dat_o[21] = wbs_ack_o;
 assign wbs_dat_o[22] = wbs_ack_o;
 assign wbs_dat_o[23] = wbs_ack_o;
 assign wbs_dat_o[24] = wbs_ack_o;
 assign wbs_dat_o[25] = wbs_ack_o;
 assign wbs_dat_o[26] = wbs_ack_o;
 assign wbs_dat_o[27] = wbs_ack_o;
 assign wbs_dat_o[28] = wbs_ack_o;
 assign wbs_dat_o[29] = wbs_ack_o;
 assign wbs_dat_o[2] = wbs_ack_o;
 assign wbs_dat_o[30] = wbs_ack_o;
 assign wbs_dat_o[31] = wbs_ack_o;
 assign wbs_dat_o[3] = wbs_ack_o;
 assign wbs_dat_o[4] = wbs_ack_o;
 assign wbs_dat_o[5] = wbs_ack_o;
 assign wbs_dat_o[6] = wbs_ack_o;
 assign wbs_dat_o[7] = wbs_ack_o;
 assign wbs_dat_o[8] = wbs_ack_o;
 assign wbs_dat_o[9] = wbs_ack_o;
endmodule
