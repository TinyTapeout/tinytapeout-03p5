magic
tech sky130A
magscale 1 2
timestamp 1685738944
<< metal1 >>
rect 281810 186260 281816 186312
rect 281868 186300 281874 186312
rect 282914 186300 282920 186312
rect 281868 186272 282920 186300
rect 281868 186260 281874 186272
rect 282914 186260 282920 186272
rect 282972 186260 282978 186312
rect 281810 184152 281816 184204
rect 281868 184192 281874 184204
rect 291838 184192 291844 184204
rect 281868 184164 291844 184192
rect 281868 184152 281874 184164
rect 291838 184152 291844 184164
rect 291896 184152 291902 184204
rect 282822 182792 282828 182844
rect 282880 182832 282886 182844
rect 288618 182832 288624 182844
rect 282880 182804 288624 182832
rect 282880 182792 282886 182804
rect 288618 182792 288624 182804
rect 288676 182832 288682 182844
rect 300854 182832 300860 182844
rect 288676 182804 300860 182832
rect 288676 182792 288682 182804
rect 300854 182792 300860 182804
rect 300912 182792 300918 182844
rect 281810 182248 281816 182300
rect 281868 182288 281874 182300
rect 285674 182288 285680 182300
rect 281868 182260 285680 182288
rect 281868 182248 281874 182260
rect 285674 182248 285680 182260
rect 285732 182248 285738 182300
rect 283558 153824 283564 153876
rect 283616 153864 283622 153876
rect 309042 153864 309048 153876
rect 283616 153836 309048 153864
rect 283616 153824 283622 153836
rect 309042 153824 309048 153836
rect 309100 153824 309106 153876
rect 309042 152464 309048 152516
rect 309100 152504 309106 152516
rect 317414 152504 317420 152516
rect 309100 152476 317420 152504
rect 309100 152464 309106 152476
rect 317414 152464 317420 152476
rect 317472 152464 317478 152516
rect 284110 72428 284116 72480
rect 284168 72468 284174 72480
rect 317414 72468 317420 72480
rect 284168 72440 317420 72468
rect 284168 72428 284174 72440
rect 317414 72428 317420 72440
rect 317472 72428 317478 72480
rect 582006 552 582012 604
rect 582064 592 582070 604
rect 583386 592 583392 604
rect 582064 564 583392 592
rect 582064 552 582070 564
rect 583386 552 583392 564
rect 583444 552 583450 604
<< via1 >>
rect 281816 186260 281868 186312
rect 282920 186260 282972 186312
rect 281816 184152 281868 184204
rect 291844 184152 291896 184204
rect 282828 182792 282880 182844
rect 288624 182792 288676 182844
rect 300860 182792 300912 182844
rect 281816 182248 281868 182300
rect 285680 182248 285732 182300
rect 283564 153824 283616 153876
rect 309048 153824 309100 153876
rect 309048 152464 309100 152516
rect 317420 152464 317472 152516
rect 284116 72428 284168 72480
rect 317420 72428 317472 72480
rect 582012 552 582064 604
rect 583392 552 583444 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 701049 8156 703520
rect 3422 701040 3478 701049
rect 3422 700975 3478 700984
rect 8114 701040 8170 701049
rect 8114 700975 8170 700984
rect 3436 254017 3464 700975
rect 24320 280809 24348 703520
rect 72988 701049 73016 703520
rect 72974 701040 73030 701049
rect 72974 700975 73030 700984
rect 89180 280945 89208 703520
rect 137848 701049 137876 703520
rect 137834 701040 137890 701049
rect 137834 700975 137890 700984
rect 154132 281081 154160 703520
rect 202800 701049 202828 703520
rect 202786 701040 202842 701049
rect 202786 700975 202842 700984
rect 154118 281072 154174 281081
rect 154118 281007 154174 281016
rect 89166 280936 89222 280945
rect 89166 280871 89222 280880
rect 24306 280800 24362 280809
rect 24306 280735 24362 280744
rect 2778 254008 2834 254017
rect 2778 253943 2834 253952
rect 3422 254008 3478 254017
rect 3422 253943 3478 253952
rect 2792 201929 2820 253943
rect 218992 214577 219020 703520
rect 267660 701049 267688 703520
rect 267646 701040 267702 701049
rect 267646 700975 267702 700984
rect 218978 214568 219034 214577
rect 218978 214503 219034 214512
rect 2778 201920 2834 201929
rect 2778 201855 2834 201864
rect 2792 188873 2820 201855
rect 283852 192545 283880 703520
rect 332520 701049 332548 703520
rect 332506 701040 332562 701049
rect 332506 700975 332562 700984
rect 348804 700505 348832 703520
rect 397472 701049 397500 703520
rect 397458 701040 397514 701049
rect 397458 700975 397514 700984
rect 292486 700496 292542 700505
rect 292486 700431 292542 700440
rect 348790 700496 348846 700505
rect 348790 700431 348846 700440
rect 289726 697504 289782 697513
rect 289726 697439 289782 697448
rect 283838 192536 283894 192545
rect 283838 192471 283894 192480
rect 287058 191992 287114 192001
rect 287058 191927 287114 191936
rect 281814 191856 281870 191865
rect 281814 191791 281870 191800
rect 9862 190360 9918 190369
rect 9862 190295 9918 190304
rect 2778 188864 2834 188873
rect 2778 188799 2834 188808
rect 2792 149841 2820 188799
rect 2778 149832 2834 149841
rect 2778 149767 2834 149776
rect 2792 97617 2820 149767
rect 2778 97608 2834 97617
rect 2778 97543 2834 97552
rect 2792 84697 2820 97543
rect 2778 84688 2834 84697
rect 2778 84623 2834 84632
rect 2792 58585 2820 84623
rect 2778 58576 2834 58585
rect 2778 58511 2834 58520
rect 2792 19417 2820 58511
rect 9876 20505 9904 190295
rect 281828 187921 281856 191791
rect 281906 190768 281962 190777
rect 281906 190703 281962 190712
rect 281814 187912 281870 187921
rect 281814 187847 281870 187856
rect 281814 186824 281870 186833
rect 281814 186759 281870 186768
rect 281828 186318 281856 186759
rect 281920 186697 281948 190703
rect 284298 189408 284354 189417
rect 284298 189343 284354 189352
rect 284312 187513 284340 189343
rect 284298 187504 284354 187513
rect 284298 187439 284354 187448
rect 285586 186824 285642 186833
rect 285586 186759 285642 186768
rect 281906 186688 281962 186697
rect 281906 186623 281962 186632
rect 281816 186312 281868 186318
rect 281816 186254 281868 186260
rect 282920 186312 282972 186318
rect 282920 186254 282972 186260
rect 282932 184793 282960 186254
rect 282918 184784 282974 184793
rect 282918 184719 282974 184728
rect 284206 184784 284262 184793
rect 284206 184719 284262 184728
rect 281814 184240 281870 184249
rect 281814 184175 281816 184184
rect 281868 184175 281870 184184
rect 281816 184146 281868 184152
rect 284114 183560 284170 183569
rect 284114 183495 284170 183504
rect 284128 183297 284156 183495
rect 282826 183288 282882 183297
rect 282826 183223 282882 183232
rect 284114 183288 284170 183297
rect 284114 183223 284170 183232
rect 282840 182850 282868 183223
rect 282828 182844 282880 182850
rect 282828 182786 282880 182792
rect 281814 182608 281870 182617
rect 281814 182543 281870 182552
rect 281828 182306 281856 182543
rect 281816 182300 281868 182306
rect 281816 182242 281868 182248
rect 281906 181928 281962 181937
rect 281906 181863 281962 181872
rect 281814 181384 281870 181393
rect 281552 181342 281814 181370
rect 281552 179466 281580 181342
rect 281814 181319 281870 181328
rect 281630 180024 281686 180033
rect 281630 179959 281686 179968
rect 281460 179438 281580 179466
rect 281460 175137 281488 179438
rect 281644 176633 281672 179959
rect 281920 179353 281948 181863
rect 281906 179344 281962 179353
rect 281906 179279 281962 179288
rect 282826 179072 282882 179081
rect 282826 179007 282882 179016
rect 281630 176624 281686 176633
rect 281630 176559 281686 176568
rect 281446 175128 281502 175137
rect 281446 175063 281502 175072
rect 282840 71369 282868 179007
rect 284220 177449 284248 184719
rect 285600 180033 285628 186759
rect 287072 184793 287100 191927
rect 288346 184920 288402 184929
rect 288346 184855 288402 184864
rect 287058 184784 287114 184793
rect 287058 184719 287114 184728
rect 285680 182300 285732 182306
rect 285680 182242 285732 182248
rect 285586 180024 285642 180033
rect 285586 179959 285642 179968
rect 285692 179217 285720 182242
rect 288360 180169 288388 184855
rect 288624 182844 288676 182850
rect 288624 182786 288676 182792
rect 288636 182209 288664 182786
rect 288622 182200 288678 182209
rect 288622 182135 288678 182144
rect 289740 180794 289768 697439
rect 290462 192536 290518 192545
rect 290462 192471 290518 192480
rect 289648 180766 289768 180794
rect 288346 180160 288402 180169
rect 288346 180095 288402 180104
rect 285678 179208 285734 179217
rect 285678 179143 285734 179152
rect 289648 177585 289676 180766
rect 289634 177576 289690 177585
rect 289634 177511 289690 177520
rect 284206 177440 284262 177449
rect 284206 177375 284262 177384
rect 283562 175128 283618 175137
rect 283562 175063 283618 175072
rect 283576 153882 283604 175063
rect 283564 153876 283616 153882
rect 283564 153818 283616 153824
rect 284116 72480 284168 72486
rect 284116 72422 284168 72428
rect 282826 71360 282882 71369
rect 282826 71295 282882 71304
rect 130566 71088 130622 71097
rect 130566 71023 130622 71032
rect 126978 69048 127034 69057
rect 126978 68983 127034 68992
rect 9862 20496 9918 20505
rect 9862 20431 9918 20440
rect 2778 19408 2834 19417
rect 2778 19343 2834 19352
rect 2792 6497 2820 19343
rect 2778 6488 2834 6497
rect 2778 6423 2834 6432
rect 2792 2825 2820 6423
rect 2778 2816 2834 2825
rect 9954 2816 10010 2825
rect 2834 2774 2912 2802
rect 2778 2751 2834 2760
rect 2884 480 2912 2774
rect 9954 2751 10010 2760
rect 14738 2816 14794 2825
rect 14738 2751 14794 2760
rect 19430 2816 19486 2825
rect 19430 2751 19486 2760
rect 24214 2816 24270 2825
rect 24214 2751 24270 2760
rect 28906 2816 28962 2825
rect 28906 2751 28962 2760
rect 32402 2816 32458 2825
rect 32402 2751 32458 2760
rect 35990 2816 36046 2825
rect 35990 2751 36046 2760
rect 39578 2816 39634 2825
rect 39578 2751 39634 2760
rect 43074 2816 43130 2825
rect 43074 2751 43130 2760
rect 46662 2816 46718 2825
rect 46662 2751 46718 2760
rect 50158 2816 50214 2825
rect 50158 2751 50214 2760
rect 53746 2816 53802 2825
rect 53746 2751 53802 2760
rect 57242 2816 57298 2825
rect 57242 2751 57298 2760
rect 60830 2816 60886 2825
rect 60830 2751 60886 2760
rect 64326 2816 64382 2825
rect 64326 2751 64382 2760
rect 67914 2816 67970 2825
rect 67914 2751 67970 2760
rect 71502 2816 71558 2825
rect 71502 2751 71558 2760
rect 74998 2816 75054 2825
rect 74998 2751 75054 2760
rect 78586 2816 78642 2825
rect 78586 2751 78642 2760
rect 82082 2816 82138 2825
rect 82082 2751 82138 2760
rect 85670 2816 85726 2825
rect 85670 2751 85726 2760
rect 89166 2816 89222 2825
rect 89166 2751 89222 2760
rect 92754 2816 92810 2825
rect 92754 2751 92810 2760
rect 96250 2816 96306 2825
rect 96250 2751 96306 2760
rect 99838 2816 99894 2825
rect 99838 2751 99894 2760
rect 103334 2816 103390 2825
rect 103334 2751 103390 2760
rect 106922 2816 106978 2825
rect 106922 2751 106978 2760
rect 110510 2816 110566 2825
rect 110510 2751 110566 2760
rect 114006 2816 114062 2825
rect 114006 2751 114062 2760
rect 117594 2816 117650 2825
rect 117594 2751 117650 2760
rect 121090 2816 121146 2825
rect 121090 2751 121146 2760
rect 124678 2816 124734 2825
rect 124678 2751 124734 2760
rect 9968 480 9996 2751
rect 14752 480 14780 2751
rect 19444 480 19472 2751
rect 24228 480 24256 2751
rect 28920 480 28948 2751
rect 32416 480 32444 2751
rect 36004 480 36032 2751
rect 39592 480 39620 2751
rect 43088 480 43116 2751
rect 46676 480 46704 2751
rect 50172 480 50200 2751
rect 53760 480 53788 2751
rect 57256 480 57284 2751
rect 60844 480 60872 2751
rect 64340 480 64368 2751
rect 67928 480 67956 2751
rect 71516 480 71544 2751
rect 75012 480 75040 2751
rect 78600 480 78628 2751
rect 82096 480 82124 2751
rect 85684 480 85712 2751
rect 89180 480 89208 2751
rect 92768 480 92796 2751
rect 96264 480 96292 2751
rect 99852 480 99880 2751
rect 103348 480 103376 2751
rect 106936 480 106964 2751
rect 110524 480 110552 2751
rect 114020 480 114048 2751
rect 117608 480 117636 2751
rect 121104 480 121132 2751
rect 124692 480 124720 2751
rect 126992 480 127020 68983
rect 130580 480 130608 71023
rect 134154 69184 134210 69193
rect 134154 69119 134210 69128
rect 134168 480 134196 69119
rect 284128 68785 284156 72422
rect 284114 68776 284170 68785
rect 284114 68711 284170 68720
rect 290476 68377 290504 192471
rect 291842 186824 291898 186833
rect 291842 186759 291898 186768
rect 291856 186425 291884 186759
rect 291842 186416 291898 186425
rect 291842 186351 291898 186360
rect 291844 184204 291896 184210
rect 291844 184146 291896 184152
rect 291856 183841 291884 184146
rect 291842 183832 291898 183841
rect 291842 183767 291898 183776
rect 292500 156777 292528 700431
rect 413664 700369 413692 703520
rect 462332 701049 462360 703520
rect 462318 701040 462374 701049
rect 462318 700975 462374 700984
rect 413650 700360 413706 700369
rect 413650 700295 413706 700304
rect 478524 697513 478552 703520
rect 527192 701049 527220 703520
rect 543476 701049 543504 703520
rect 527178 701040 527234 701049
rect 527178 700975 527234 700984
rect 543462 701040 543518 701049
rect 543462 700975 543518 700984
rect 543476 697513 543504 700975
rect 559668 700369 559696 703520
rect 559654 700360 559710 700369
rect 559654 700295 559710 700304
rect 582378 700360 582434 700369
rect 582378 700295 582434 700304
rect 478510 697504 478566 697513
rect 478510 697439 478566 697448
rect 543462 697504 543518 697513
rect 543462 697439 543518 697448
rect 580906 697232 580962 697241
rect 580906 697167 580962 697176
rect 580920 683913 580948 697167
rect 580906 683904 580962 683913
rect 580906 683839 580962 683848
rect 580920 644065 580948 683839
rect 580906 644056 580962 644065
rect 580906 643991 580962 644000
rect 580920 630873 580948 643991
rect 580906 630864 580962 630873
rect 580906 630799 580962 630808
rect 580920 591025 580948 630799
rect 580906 591016 580962 591025
rect 580906 590951 580962 590960
rect 580920 577697 580948 590951
rect 580906 577688 580962 577697
rect 580906 577623 580962 577632
rect 580920 537849 580948 577623
rect 580906 537840 580962 537849
rect 580906 537775 580962 537784
rect 580920 524521 580948 537775
rect 580906 524512 580962 524521
rect 580906 524447 580962 524456
rect 580920 484673 580948 524447
rect 580906 484664 580962 484673
rect 580906 484599 580962 484608
rect 580920 471481 580948 484599
rect 580906 471472 580962 471481
rect 580906 471407 580962 471416
rect 580920 431633 580948 471407
rect 580906 431624 580962 431633
rect 580906 431559 580962 431568
rect 580920 418305 580948 431559
rect 580906 418296 580962 418305
rect 580906 418231 580962 418240
rect 580920 378457 580948 418231
rect 580906 378448 580962 378457
rect 580906 378383 580962 378392
rect 580920 365129 580948 378383
rect 580906 365120 580962 365129
rect 580906 365055 580962 365064
rect 580920 325281 580948 365055
rect 580906 325272 580962 325281
rect 580906 325207 580962 325216
rect 439134 323504 439190 323513
rect 439134 323439 439190 323448
rect 439148 319841 439176 323439
rect 439134 319832 439190 319841
rect 439134 319767 439190 319776
rect 580920 312089 580948 325207
rect 580906 312080 580962 312089
rect 580906 312015 580962 312024
rect 580920 272241 580948 312015
rect 580906 272232 580962 272241
rect 580906 272167 580962 272176
rect 580920 259457 580948 272167
rect 580906 259448 580962 259457
rect 580906 259383 580962 259392
rect 300766 247072 300822 247081
rect 300766 247007 300822 247016
rect 300780 220969 300808 247007
rect 580906 232384 580962 232393
rect 580906 232319 580962 232328
rect 300766 220960 300822 220969
rect 300766 220895 300822 220904
rect 307758 220960 307814 220969
rect 307758 220895 307814 220904
rect 307772 212945 307800 220895
rect 327722 215792 327778 215801
rect 327722 215727 327778 215736
rect 327736 212945 327764 215727
rect 307758 212936 307814 212945
rect 307758 212871 307814 212880
rect 327722 212936 327778 212945
rect 327722 212871 327778 212880
rect 580920 192545 580948 232319
rect 580906 192536 580962 192545
rect 580906 192471 580962 192480
rect 298098 191992 298154 192001
rect 298098 191927 298154 191936
rect 297546 189136 297602 189145
rect 297546 189071 297602 189080
rect 295982 187776 296038 187785
rect 295982 187711 296038 187720
rect 292486 156768 292542 156777
rect 292486 156703 292542 156712
rect 295996 71097 296024 187711
rect 297560 186153 297588 189071
rect 298112 186833 298140 191927
rect 300490 190632 300546 190641
rect 300490 190567 300546 190576
rect 300504 189281 300532 190567
rect 302330 190496 302386 190505
rect 302330 190431 302386 190440
rect 300950 189544 301006 189553
rect 300950 189479 301006 189488
rect 300490 189272 300546 189281
rect 300490 189207 300546 189216
rect 298190 186960 298246 186969
rect 298190 186895 298246 186904
rect 298098 186824 298154 186833
rect 298098 186759 298154 186768
rect 297546 186144 297602 186153
rect 297546 186079 297602 186088
rect 296626 180432 296682 180441
rect 296626 180367 296682 180376
rect 296640 176633 296668 180367
rect 296626 176624 296682 176633
rect 296626 176559 296682 176568
rect 296626 167104 296682 167113
rect 296626 167039 296682 167048
rect 296640 161537 296668 167039
rect 296626 161528 296682 161537
rect 296626 161463 296682 161472
rect 296626 161392 296682 161401
rect 296626 161327 296682 161336
rect 296640 151881 296668 161327
rect 296626 151872 296682 151881
rect 296626 151807 296682 151816
rect 295982 71088 296038 71097
rect 295982 71023 296038 71032
rect 290462 68368 290518 68377
rect 290462 68303 290518 68312
rect 273902 67960 273958 67969
rect 273902 67895 273958 67904
rect 271142 67824 271198 67833
rect 271142 67759 271198 67768
rect 151818 67688 151874 67697
rect 151818 67623 151874 67632
rect 137650 65920 137706 65929
rect 137650 65855 137706 65864
rect 137664 480 137692 65855
rect 148322 65784 148378 65793
rect 148322 65719 148378 65728
rect 144734 64288 144790 64297
rect 144734 64223 144790 64232
rect 141238 64152 141294 64161
rect 141238 64087 141294 64096
rect 141252 480 141280 64087
rect 144748 480 144776 64223
rect 148336 480 148364 65719
rect 151832 480 151860 67623
rect 158902 66328 158958 66337
rect 158902 66263 158958 66272
rect 155406 62792 155462 62801
rect 155406 62727 155462 62736
rect 155420 480 155448 62727
rect 158916 480 158944 66263
rect 271156 64161 271184 67759
rect 273916 64297 273944 67895
rect 297560 67561 297588 186079
rect 298204 180794 298232 186895
rect 300766 184648 300822 184657
rect 300766 184583 300822 184592
rect 299570 184240 299626 184249
rect 299570 184175 299626 184184
rect 299584 183841 299612 184175
rect 299570 183832 299626 183841
rect 299570 183767 299626 183776
rect 298112 180766 298232 180794
rect 298112 67697 298140 180766
rect 300780 179489 300808 184583
rect 300858 183288 300914 183297
rect 300858 183223 300914 183232
rect 300872 182850 300900 183223
rect 300860 182844 300912 182850
rect 300860 182786 300912 182792
rect 300964 181393 300992 189479
rect 302238 189272 302294 189281
rect 302238 189207 302294 189216
rect 302252 187377 302280 189207
rect 302238 187368 302294 187377
rect 302238 187303 302294 187312
rect 302252 186314 302280 187303
rect 302344 186697 302372 190431
rect 302330 186688 302386 186697
rect 302330 186623 302386 186632
rect 302252 186286 302372 186314
rect 302238 181928 302294 181937
rect 302238 181863 302294 181872
rect 300950 181384 301006 181393
rect 300950 181319 301006 181328
rect 302252 179738 302280 181863
rect 302344 180794 302372 186286
rect 302344 180766 302648 180794
rect 302252 179710 302372 179738
rect 302238 179616 302294 179625
rect 302238 179551 302294 179560
rect 300766 179480 300822 179489
rect 300766 179415 300822 179424
rect 301502 179480 301558 179489
rect 301502 179415 301558 179424
rect 301516 156641 301544 179415
rect 301502 156632 301558 156641
rect 301502 156567 301558 156576
rect 302252 69034 302280 179551
rect 302344 179353 302372 179710
rect 302330 179344 302386 179353
rect 302330 179279 302386 179288
rect 302344 178945 302372 179279
rect 302620 179217 302648 180766
rect 580920 179217 580948 192471
rect 302606 179208 302662 179217
rect 302606 179143 302662 179152
rect 580906 179208 580962 179217
rect 580906 179143 580962 179152
rect 302330 178936 302386 178945
rect 302330 178871 302386 178880
rect 311898 157856 311954 157865
rect 311898 157791 311954 157800
rect 306378 157312 306434 157321
rect 306378 157247 306434 157256
rect 303618 156632 303674 156641
rect 303618 156567 303674 156576
rect 302160 69006 302280 69034
rect 302160 68785 302188 69006
rect 302146 68776 302202 68785
rect 302146 68711 302202 68720
rect 303632 68513 303660 156567
rect 304998 71360 305054 71369
rect 304998 71295 305054 71304
rect 303618 68504 303674 68513
rect 303618 68439 303674 68448
rect 298098 67688 298154 67697
rect 298098 67623 298154 67632
rect 305012 67561 305040 71295
rect 306392 68649 306420 157247
rect 309138 157040 309194 157049
rect 309138 156975 309194 156984
rect 309048 153876 309100 153882
rect 309048 153818 309100 153824
rect 309060 152522 309088 153818
rect 309048 152516 309100 152522
rect 309048 152458 309100 152464
rect 306378 68640 306434 68649
rect 306378 68575 306434 68584
rect 297546 67552 297602 67561
rect 297546 67487 297602 67496
rect 304998 67552 305054 67561
rect 304998 67487 305054 67496
rect 309152 67017 309180 156975
rect 311912 68921 311940 157791
rect 317420 152516 317472 152522
rect 317420 152458 317472 152464
rect 317432 72486 317460 152458
rect 317420 72480 317472 72486
rect 317420 72422 317472 72428
rect 311898 68912 311954 68921
rect 311898 68847 311954 68856
rect 309138 67008 309194 67017
rect 309138 66943 309194 66952
rect 279882 66600 279938 66609
rect 279882 66535 279938 66544
rect 279896 65793 279924 66535
rect 279882 65784 279938 65793
rect 279882 65719 279938 65728
rect 273902 64288 273958 64297
rect 273902 64223 273958 64232
rect 271142 64152 271198 64161
rect 271142 64087 271198 64096
rect 273902 44840 273958 44849
rect 273902 44775 273958 44784
rect 273916 22001 273944 44775
rect 273902 21992 273958 22001
rect 273902 21927 273958 21936
rect 278686 21992 278742 22001
rect 278686 21927 278742 21936
rect 278700 20505 278728 21927
rect 278686 20496 278742 20505
rect 278686 20431 278742 20440
rect 277306 19544 277362 19553
rect 277306 19479 277362 19488
rect 277320 19145 277348 19479
rect 278042 19408 278098 19417
rect 278042 19343 278098 19352
rect 277306 19136 277362 19145
rect 277306 19071 277362 19080
rect 278056 2825 278084 19343
rect 579802 3496 579858 3505
rect 579802 3431 579858 3440
rect 570326 3360 570382 3369
rect 570326 3295 570382 3304
rect 573914 3360 573970 3369
rect 573914 3295 573970 3304
rect 577410 3360 577466 3369
rect 577410 3295 577466 3304
rect 162490 2816 162546 2825
rect 162490 2751 162546 2760
rect 166078 2816 166134 2825
rect 166078 2751 166134 2760
rect 169574 2816 169630 2825
rect 169574 2751 169630 2760
rect 173162 2816 173218 2825
rect 173162 2751 173218 2760
rect 176658 2816 176714 2825
rect 176658 2751 176714 2760
rect 180246 2816 180302 2825
rect 180246 2751 180302 2760
rect 183742 2816 183798 2825
rect 183742 2751 183798 2760
rect 187330 2816 187386 2825
rect 187330 2751 187386 2760
rect 190826 2816 190882 2825
rect 190826 2751 190882 2760
rect 194414 2816 194470 2825
rect 194414 2751 194470 2760
rect 197910 2816 197966 2825
rect 197910 2751 197966 2760
rect 201498 2816 201554 2825
rect 201498 2751 201554 2760
rect 205086 2816 205142 2825
rect 205086 2751 205142 2760
rect 208582 2816 208638 2825
rect 208582 2751 208638 2760
rect 212170 2816 212226 2825
rect 212170 2751 212226 2760
rect 215666 2816 215722 2825
rect 215666 2751 215722 2760
rect 219254 2816 219310 2825
rect 219254 2751 219310 2760
rect 222750 2816 222806 2825
rect 222750 2751 222806 2760
rect 226338 2816 226394 2825
rect 226338 2751 226394 2760
rect 229834 2816 229890 2825
rect 229834 2751 229890 2760
rect 233422 2816 233478 2825
rect 233422 2751 233478 2760
rect 237010 2816 237066 2825
rect 237010 2751 237066 2760
rect 240506 2816 240562 2825
rect 240506 2751 240562 2760
rect 244094 2816 244150 2825
rect 244094 2751 244150 2760
rect 247590 2816 247646 2825
rect 247590 2751 247646 2760
rect 251178 2816 251234 2825
rect 251178 2751 251234 2760
rect 254674 2816 254730 2825
rect 254674 2751 254730 2760
rect 258262 2816 258318 2825
rect 258262 2751 258318 2760
rect 261758 2816 261814 2825
rect 261758 2751 261814 2760
rect 265346 2816 265402 2825
rect 265346 2751 265402 2760
rect 268842 2816 268898 2825
rect 268842 2751 268898 2760
rect 272430 2816 272486 2825
rect 272430 2751 272486 2760
rect 276018 2816 276074 2825
rect 276018 2751 276074 2760
rect 278042 2816 278098 2825
rect 278042 2751 278098 2760
rect 279514 2816 279570 2825
rect 279514 2751 279570 2760
rect 283102 2816 283158 2825
rect 283102 2751 283158 2760
rect 286598 2816 286654 2825
rect 286598 2751 286654 2760
rect 290186 2816 290242 2825
rect 290186 2751 290242 2760
rect 293682 2816 293738 2825
rect 293682 2751 293738 2760
rect 297270 2816 297326 2825
rect 297270 2751 297326 2760
rect 300766 2816 300822 2825
rect 300766 2751 300822 2760
rect 304354 2816 304410 2825
rect 304354 2751 304410 2760
rect 307942 2816 307998 2825
rect 307942 2751 307998 2760
rect 311438 2816 311494 2825
rect 311438 2751 311494 2760
rect 315026 2816 315082 2825
rect 315026 2751 315082 2760
rect 318522 2816 318578 2825
rect 318522 2751 318578 2760
rect 322110 2816 322166 2825
rect 322110 2751 322166 2760
rect 325606 2816 325662 2825
rect 325606 2751 325662 2760
rect 329194 2816 329250 2825
rect 329194 2751 329250 2760
rect 332690 2816 332746 2825
rect 332690 2751 332746 2760
rect 336278 2816 336334 2825
rect 336278 2751 336334 2760
rect 339866 2816 339922 2825
rect 339866 2751 339922 2760
rect 343362 2816 343418 2825
rect 343362 2751 343418 2760
rect 346950 2816 347006 2825
rect 346950 2751 347006 2760
rect 350446 2816 350502 2825
rect 350446 2751 350502 2760
rect 354034 2816 354090 2825
rect 354034 2751 354090 2760
rect 357530 2816 357586 2825
rect 357530 2751 357586 2760
rect 361118 2816 361174 2825
rect 361118 2751 361174 2760
rect 364614 2816 364670 2825
rect 364614 2751 364670 2760
rect 368202 2816 368258 2825
rect 368202 2751 368258 2760
rect 371698 2816 371754 2825
rect 371698 2751 371754 2760
rect 375286 2816 375342 2825
rect 375286 2751 375342 2760
rect 378874 2816 378930 2825
rect 378874 2751 378930 2760
rect 382370 2816 382426 2825
rect 382370 2751 382426 2760
rect 385958 2816 386014 2825
rect 385958 2751 386014 2760
rect 389454 2816 389510 2825
rect 389454 2751 389510 2760
rect 393042 2816 393098 2825
rect 393042 2751 393098 2760
rect 396538 2816 396594 2825
rect 396538 2751 396594 2760
rect 400126 2816 400182 2825
rect 400126 2751 400182 2760
rect 403622 2816 403678 2825
rect 403622 2751 403678 2760
rect 407210 2816 407266 2825
rect 407210 2751 407266 2760
rect 410798 2816 410854 2825
rect 410798 2751 410854 2760
rect 414294 2816 414350 2825
rect 414294 2751 414350 2760
rect 417882 2816 417938 2825
rect 417882 2751 417938 2760
rect 421378 2816 421434 2825
rect 421378 2751 421434 2760
rect 424966 2816 425022 2825
rect 424966 2751 425022 2760
rect 428462 2816 428518 2825
rect 428462 2751 428518 2760
rect 432050 2816 432106 2825
rect 432050 2751 432106 2760
rect 435546 2816 435602 2825
rect 435546 2751 435602 2760
rect 439134 2816 439190 2825
rect 439134 2751 439190 2760
rect 442630 2816 442686 2825
rect 442630 2751 442686 2760
rect 446218 2816 446274 2825
rect 446218 2751 446274 2760
rect 449806 2816 449862 2825
rect 449806 2751 449862 2760
rect 453302 2816 453358 2825
rect 453302 2751 453358 2760
rect 456890 2816 456946 2825
rect 456890 2751 456946 2760
rect 460386 2816 460442 2825
rect 460386 2751 460442 2760
rect 463974 2816 464030 2825
rect 463974 2751 464030 2760
rect 467470 2816 467526 2825
rect 467470 2751 467526 2760
rect 471058 2816 471114 2825
rect 471058 2751 471114 2760
rect 474554 2816 474610 2825
rect 474554 2751 474610 2760
rect 478142 2816 478198 2825
rect 478142 2751 478198 2760
rect 481730 2816 481786 2825
rect 481730 2751 481786 2760
rect 485226 2816 485282 2825
rect 485226 2751 485282 2760
rect 488814 2816 488870 2825
rect 488814 2751 488870 2760
rect 492310 2816 492366 2825
rect 492310 2751 492366 2760
rect 495898 2816 495954 2825
rect 495898 2751 495954 2760
rect 499394 2816 499450 2825
rect 499394 2751 499450 2760
rect 502982 2816 503038 2825
rect 502982 2751 503038 2760
rect 506478 2816 506534 2825
rect 506478 2751 506534 2760
rect 510066 2816 510122 2825
rect 510066 2751 510122 2760
rect 513562 2816 513618 2825
rect 513562 2751 513618 2760
rect 517150 2816 517206 2825
rect 517150 2751 517206 2760
rect 520738 2816 520794 2825
rect 520738 2751 520794 2760
rect 524234 2816 524290 2825
rect 524234 2751 524290 2760
rect 527822 2816 527878 2825
rect 527822 2751 527878 2760
rect 531318 2816 531374 2825
rect 531318 2751 531374 2760
rect 534906 2816 534962 2825
rect 534906 2751 534962 2760
rect 538402 2816 538458 2825
rect 538402 2751 538458 2760
rect 541990 2816 542046 2825
rect 541990 2751 542046 2760
rect 545486 2816 545542 2825
rect 545486 2751 545542 2760
rect 549074 2816 549130 2825
rect 549074 2751 549130 2760
rect 552662 2816 552718 2825
rect 552662 2751 552718 2760
rect 556158 2816 556214 2825
rect 556158 2751 556214 2760
rect 559746 2816 559802 2825
rect 559746 2751 559802 2760
rect 563242 2816 563298 2825
rect 563242 2751 563298 2760
rect 566830 2816 566886 2825
rect 566830 2751 566886 2760
rect 162504 480 162532 2751
rect 166092 480 166120 2751
rect 169588 480 169616 2751
rect 173176 480 173204 2751
rect 176672 480 176700 2751
rect 180260 480 180288 2751
rect 183756 480 183784 2751
rect 187344 480 187372 2751
rect 190840 480 190868 2751
rect 194428 480 194456 2751
rect 197924 480 197952 2751
rect 201512 480 201540 2751
rect 205100 480 205128 2751
rect 208596 480 208624 2751
rect 212184 480 212212 2751
rect 215680 480 215708 2751
rect 219268 480 219296 2751
rect 222764 480 222792 2751
rect 226352 480 226380 2751
rect 229848 480 229876 2751
rect 233436 480 233464 2751
rect 237024 480 237052 2751
rect 240520 480 240548 2751
rect 244108 480 244136 2751
rect 247604 480 247632 2751
rect 251192 480 251220 2751
rect 254688 480 254716 2751
rect 258276 480 258304 2751
rect 261772 480 261800 2751
rect 265360 480 265388 2751
rect 268856 480 268884 2751
rect 272444 480 272472 2751
rect 276032 480 276060 2751
rect 279528 480 279556 2751
rect 283116 480 283144 2751
rect 286612 480 286640 2751
rect 290200 480 290228 2751
rect 293696 480 293724 2751
rect 297284 480 297312 2751
rect 300780 480 300808 2751
rect 304368 480 304396 2751
rect 307956 480 307984 2751
rect 311452 480 311480 2751
rect 315040 480 315068 2751
rect 318536 480 318564 2751
rect 322124 480 322152 2751
rect 325620 480 325648 2751
rect 329208 480 329236 2751
rect 332704 480 332732 2751
rect 336292 480 336320 2751
rect 339880 480 339908 2751
rect 343376 480 343404 2751
rect 346964 480 346992 2751
rect 350460 480 350488 2751
rect 354048 480 354076 2751
rect 357544 480 357572 2751
rect 361132 480 361160 2751
rect 364628 480 364656 2751
rect 368216 480 368244 2751
rect 371712 480 371740 2751
rect 375300 480 375328 2751
rect 378888 480 378916 2751
rect 382384 480 382412 2751
rect 385972 480 386000 2751
rect 389468 480 389496 2751
rect 393056 480 393084 2751
rect 396552 480 396580 2751
rect 400140 480 400168 2751
rect 403636 480 403664 2751
rect 407224 480 407252 2751
rect 410812 480 410840 2751
rect 414308 480 414336 2751
rect 417896 480 417924 2751
rect 421392 480 421420 2751
rect 424980 480 425008 2751
rect 428476 480 428504 2751
rect 432064 480 432092 2751
rect 435560 480 435588 2751
rect 439148 480 439176 2751
rect 442644 480 442672 2751
rect 446232 480 446260 2751
rect 449820 480 449848 2751
rect 453316 480 453344 2751
rect 456904 480 456932 2751
rect 460400 480 460428 2751
rect 463988 480 464016 2751
rect 467484 480 467512 2751
rect 471072 480 471100 2751
rect 474568 480 474596 2751
rect 478156 480 478184 2751
rect 481744 480 481772 2751
rect 485240 480 485268 2751
rect 488828 480 488856 2751
rect 492324 480 492352 2751
rect 495912 480 495940 2751
rect 499408 480 499436 2751
rect 502996 480 503024 2751
rect 506492 480 506520 2751
rect 510080 480 510108 2751
rect 513576 480 513604 2751
rect 517164 480 517192 2751
rect 520752 480 520780 2751
rect 524248 480 524276 2751
rect 527836 480 527864 2751
rect 531332 480 531360 2751
rect 534920 480 534948 2751
rect 538416 480 538444 2751
rect 542004 480 542032 2751
rect 545500 480 545528 2751
rect 549088 480 549116 2751
rect 552676 480 552704 2751
rect 556172 480 556200 2751
rect 559760 480 559788 2751
rect 563256 480 563284 2751
rect 566844 480 566872 2751
rect 570340 480 570368 3295
rect 573928 480 573956 3295
rect 577424 480 577452 3295
rect 579816 480 579844 3431
rect 580920 3369 580948 179143
rect 582392 68241 582420 700295
rect 582378 68232 582434 68241
rect 582378 68167 582434 68176
rect 580906 3360 580962 3369
rect 580962 3318 581040 3346
rect 580906 3295 580962 3304
rect 581012 626 581040 3318
rect 581012 598 581224 626
rect 581012 480 581040 598
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 581196 354 581224 598
rect 582012 604 582064 610
rect 582012 546 582064 552
rect 583392 604 583444 610
rect 583392 546 583444 552
rect 581196 326 581776 354
rect 581748 218 581776 326
rect 582024 218 582052 546
rect 583404 480 583432 546
rect 582166 218 582278 480
rect 581748 190 582278 218
rect 582166 -960 582278 190
rect 583362 -960 583474 480
<< via2 >>
rect 3422 700984 3478 701040
rect 8114 700984 8170 701040
rect 72974 700984 73030 701040
rect 137834 700984 137890 701040
rect 202786 700984 202842 701040
rect 154118 281016 154174 281072
rect 89166 280880 89222 280936
rect 24306 280744 24362 280800
rect 2778 253952 2834 254008
rect 3422 253952 3478 254008
rect 267646 700984 267702 701040
rect 218978 214512 219034 214568
rect 2778 201864 2834 201920
rect 332506 700984 332562 701040
rect 397458 700984 397514 701040
rect 292486 700440 292542 700496
rect 348790 700440 348846 700496
rect 289726 697448 289782 697504
rect 283838 192480 283894 192536
rect 287058 191936 287114 191992
rect 281814 191800 281870 191856
rect 9862 190304 9918 190360
rect 2778 188808 2834 188864
rect 2778 149776 2834 149832
rect 2778 97552 2834 97608
rect 2778 84632 2834 84688
rect 2778 58520 2834 58576
rect 281906 190712 281962 190768
rect 281814 187856 281870 187912
rect 281814 186768 281870 186824
rect 284298 189352 284354 189408
rect 284298 187448 284354 187504
rect 285586 186768 285642 186824
rect 281906 186632 281962 186688
rect 282918 184728 282974 184784
rect 284206 184728 284262 184784
rect 281814 184204 281870 184240
rect 281814 184184 281816 184204
rect 281816 184184 281868 184204
rect 281868 184184 281870 184204
rect 284114 183504 284170 183560
rect 282826 183232 282882 183288
rect 284114 183232 284170 183288
rect 281814 182552 281870 182608
rect 281906 181872 281962 181928
rect 281814 181328 281870 181384
rect 281630 179968 281686 180024
rect 281906 179288 281962 179344
rect 282826 179016 282882 179072
rect 281630 176568 281686 176624
rect 281446 175072 281502 175128
rect 288346 184864 288402 184920
rect 287058 184728 287114 184784
rect 285586 179968 285642 180024
rect 288622 182144 288678 182200
rect 290462 192480 290518 192536
rect 288346 180104 288402 180160
rect 285678 179152 285734 179208
rect 289634 177520 289690 177576
rect 284206 177384 284262 177440
rect 283562 175072 283618 175128
rect 282826 71304 282882 71360
rect 130566 71032 130622 71088
rect 126978 68992 127034 69048
rect 9862 20440 9918 20496
rect 2778 19352 2834 19408
rect 2778 6432 2834 6488
rect 2778 2760 2834 2816
rect 9954 2760 10010 2816
rect 14738 2760 14794 2816
rect 19430 2760 19486 2816
rect 24214 2760 24270 2816
rect 28906 2760 28962 2816
rect 32402 2760 32458 2816
rect 35990 2760 36046 2816
rect 39578 2760 39634 2816
rect 43074 2760 43130 2816
rect 46662 2760 46718 2816
rect 50158 2760 50214 2816
rect 53746 2760 53802 2816
rect 57242 2760 57298 2816
rect 60830 2760 60886 2816
rect 64326 2760 64382 2816
rect 67914 2760 67970 2816
rect 71502 2760 71558 2816
rect 74998 2760 75054 2816
rect 78586 2760 78642 2816
rect 82082 2760 82138 2816
rect 85670 2760 85726 2816
rect 89166 2760 89222 2816
rect 92754 2760 92810 2816
rect 96250 2760 96306 2816
rect 99838 2760 99894 2816
rect 103334 2760 103390 2816
rect 106922 2760 106978 2816
rect 110510 2760 110566 2816
rect 114006 2760 114062 2816
rect 117594 2760 117650 2816
rect 121090 2760 121146 2816
rect 124678 2760 124734 2816
rect 134154 69128 134210 69184
rect 284114 68720 284170 68776
rect 291842 186768 291898 186824
rect 291842 186360 291898 186416
rect 291842 183776 291898 183832
rect 462318 700984 462374 701040
rect 413650 700304 413706 700360
rect 527178 700984 527234 701040
rect 543462 700984 543518 701040
rect 559654 700304 559710 700360
rect 582378 700304 582434 700360
rect 478510 697448 478566 697504
rect 543462 697448 543518 697504
rect 580906 697176 580962 697232
rect 580906 683848 580962 683904
rect 580906 644000 580962 644056
rect 580906 630808 580962 630864
rect 580906 590960 580962 591016
rect 580906 577632 580962 577688
rect 580906 537784 580962 537840
rect 580906 524456 580962 524512
rect 580906 484608 580962 484664
rect 580906 471416 580962 471472
rect 580906 431568 580962 431624
rect 580906 418240 580962 418296
rect 580906 378392 580962 378448
rect 580906 365064 580962 365120
rect 580906 325216 580962 325272
rect 439134 323448 439190 323504
rect 439134 319776 439190 319832
rect 580906 312024 580962 312080
rect 580906 272176 580962 272232
rect 580906 259392 580962 259448
rect 300766 247016 300822 247072
rect 580906 232328 580962 232384
rect 300766 220904 300822 220960
rect 307758 220904 307814 220960
rect 327722 215736 327778 215792
rect 307758 212880 307814 212936
rect 327722 212880 327778 212936
rect 580906 192480 580962 192536
rect 298098 191936 298154 191992
rect 297546 189080 297602 189136
rect 295982 187720 296038 187776
rect 292486 156712 292542 156768
rect 300490 190576 300546 190632
rect 302330 190440 302386 190496
rect 300950 189488 301006 189544
rect 300490 189216 300546 189272
rect 298190 186904 298246 186960
rect 298098 186768 298154 186824
rect 297546 186088 297602 186144
rect 296626 180376 296682 180432
rect 296626 176568 296682 176624
rect 296626 167048 296682 167104
rect 296626 161472 296682 161528
rect 296626 161336 296682 161392
rect 296626 151816 296682 151872
rect 295982 71032 296038 71088
rect 290462 68312 290518 68368
rect 273902 67904 273958 67960
rect 271142 67768 271198 67824
rect 151818 67632 151874 67688
rect 137650 65864 137706 65920
rect 148322 65728 148378 65784
rect 144734 64232 144790 64288
rect 141238 64096 141294 64152
rect 158902 66272 158958 66328
rect 155406 62736 155462 62792
rect 300766 184592 300822 184648
rect 299570 184184 299626 184240
rect 299570 183776 299626 183832
rect 300858 183232 300914 183288
rect 302238 189216 302294 189272
rect 302238 187312 302294 187368
rect 302330 186632 302386 186688
rect 302238 181872 302294 181928
rect 300950 181328 301006 181384
rect 302238 179560 302294 179616
rect 300766 179424 300822 179480
rect 301502 179424 301558 179480
rect 301502 156576 301558 156632
rect 302330 179288 302386 179344
rect 302606 179152 302662 179208
rect 580906 179152 580962 179208
rect 302330 178880 302386 178936
rect 311898 157800 311954 157856
rect 306378 157256 306434 157312
rect 303618 156576 303674 156632
rect 302146 68720 302202 68776
rect 304998 71304 305054 71360
rect 303618 68448 303674 68504
rect 298098 67632 298154 67688
rect 309138 156984 309194 157040
rect 306378 68584 306434 68640
rect 297546 67496 297602 67552
rect 304998 67496 305054 67552
rect 311898 68856 311954 68912
rect 309138 66952 309194 67008
rect 279882 66544 279938 66600
rect 279882 65728 279938 65784
rect 273902 64232 273958 64288
rect 271142 64096 271198 64152
rect 273902 44784 273958 44840
rect 273902 21936 273958 21992
rect 278686 21936 278742 21992
rect 278686 20440 278742 20496
rect 277306 19488 277362 19544
rect 278042 19352 278098 19408
rect 277306 19080 277362 19136
rect 579802 3440 579858 3496
rect 570326 3304 570382 3360
rect 573914 3304 573970 3360
rect 577410 3304 577466 3360
rect 162490 2760 162546 2816
rect 166078 2760 166134 2816
rect 169574 2760 169630 2816
rect 173162 2760 173218 2816
rect 176658 2760 176714 2816
rect 180246 2760 180302 2816
rect 183742 2760 183798 2816
rect 187330 2760 187386 2816
rect 190826 2760 190882 2816
rect 194414 2760 194470 2816
rect 197910 2760 197966 2816
rect 201498 2760 201554 2816
rect 205086 2760 205142 2816
rect 208582 2760 208638 2816
rect 212170 2760 212226 2816
rect 215666 2760 215722 2816
rect 219254 2760 219310 2816
rect 222750 2760 222806 2816
rect 226338 2760 226394 2816
rect 229834 2760 229890 2816
rect 233422 2760 233478 2816
rect 237010 2760 237066 2816
rect 240506 2760 240562 2816
rect 244094 2760 244150 2816
rect 247590 2760 247646 2816
rect 251178 2760 251234 2816
rect 254674 2760 254730 2816
rect 258262 2760 258318 2816
rect 261758 2760 261814 2816
rect 265346 2760 265402 2816
rect 268842 2760 268898 2816
rect 272430 2760 272486 2816
rect 276018 2760 276074 2816
rect 278042 2760 278098 2816
rect 279514 2760 279570 2816
rect 283102 2760 283158 2816
rect 286598 2760 286654 2816
rect 290186 2760 290242 2816
rect 293682 2760 293738 2816
rect 297270 2760 297326 2816
rect 300766 2760 300822 2816
rect 304354 2760 304410 2816
rect 307942 2760 307998 2816
rect 311438 2760 311494 2816
rect 315026 2760 315082 2816
rect 318522 2760 318578 2816
rect 322110 2760 322166 2816
rect 325606 2760 325662 2816
rect 329194 2760 329250 2816
rect 332690 2760 332746 2816
rect 336278 2760 336334 2816
rect 339866 2760 339922 2816
rect 343362 2760 343418 2816
rect 346950 2760 347006 2816
rect 350446 2760 350502 2816
rect 354034 2760 354090 2816
rect 357530 2760 357586 2816
rect 361118 2760 361174 2816
rect 364614 2760 364670 2816
rect 368202 2760 368258 2816
rect 371698 2760 371754 2816
rect 375286 2760 375342 2816
rect 378874 2760 378930 2816
rect 382370 2760 382426 2816
rect 385958 2760 386014 2816
rect 389454 2760 389510 2816
rect 393042 2760 393098 2816
rect 396538 2760 396594 2816
rect 400126 2760 400182 2816
rect 403622 2760 403678 2816
rect 407210 2760 407266 2816
rect 410798 2760 410854 2816
rect 414294 2760 414350 2816
rect 417882 2760 417938 2816
rect 421378 2760 421434 2816
rect 424966 2760 425022 2816
rect 428462 2760 428518 2816
rect 432050 2760 432106 2816
rect 435546 2760 435602 2816
rect 439134 2760 439190 2816
rect 442630 2760 442686 2816
rect 446218 2760 446274 2816
rect 449806 2760 449862 2816
rect 453302 2760 453358 2816
rect 456890 2760 456946 2816
rect 460386 2760 460442 2816
rect 463974 2760 464030 2816
rect 467470 2760 467526 2816
rect 471058 2760 471114 2816
rect 474554 2760 474610 2816
rect 478142 2760 478198 2816
rect 481730 2760 481786 2816
rect 485226 2760 485282 2816
rect 488814 2760 488870 2816
rect 492310 2760 492366 2816
rect 495898 2760 495954 2816
rect 499394 2760 499450 2816
rect 502982 2760 503038 2816
rect 506478 2760 506534 2816
rect 510066 2760 510122 2816
rect 513562 2760 513618 2816
rect 517150 2760 517206 2816
rect 520738 2760 520794 2816
rect 524234 2760 524290 2816
rect 527822 2760 527878 2816
rect 531318 2760 531374 2816
rect 534906 2760 534962 2816
rect 538402 2760 538458 2816
rect 541990 2760 542046 2816
rect 545486 2760 545542 2816
rect 549074 2760 549130 2816
rect 552662 2760 552718 2816
rect 556158 2760 556214 2816
rect 559746 2760 559802 2816
rect 563242 2760 563298 2816
rect 566830 2760 566886 2816
rect 582378 68176 582434 68232
rect 580906 3304 580962 3360
<< metal3 >>
rect 3417 701042 3483 701045
rect 8109 701042 8175 701045
rect 72969 701042 73035 701045
rect 137829 701042 137895 701045
rect 202781 701042 202847 701045
rect 267641 701042 267707 701045
rect 332501 701042 332567 701045
rect 397453 701042 397519 701045
rect 462313 701042 462379 701045
rect 3417 701040 462379 701042
rect 3417 700984 3422 701040
rect 3478 700984 8114 701040
rect 8170 700984 72974 701040
rect 73030 700984 137834 701040
rect 137890 700984 202786 701040
rect 202842 700984 267646 701040
rect 267702 700984 332506 701040
rect 332562 700984 397458 701040
rect 397514 700984 462318 701040
rect 462374 700984 462379 701040
rect 3417 700982 462379 700984
rect 3417 700979 3483 700982
rect 8109 700979 8175 700982
rect 72969 700979 73035 700982
rect 137829 700979 137895 700982
rect 202781 700979 202847 700982
rect 267641 700979 267707 700982
rect 332501 700979 332567 700982
rect 397453 700979 397519 700982
rect 462313 700979 462379 700982
rect 527173 701042 527239 701045
rect 543457 701042 543523 701045
rect 527173 701040 543523 701042
rect 527173 700984 527178 701040
rect 527234 700984 543462 701040
rect 543518 700984 543523 701040
rect 527173 700982 543523 700984
rect 527173 700979 527239 700982
rect 543457 700979 543523 700982
rect 292481 700498 292547 700501
rect 348785 700498 348851 700501
rect 292481 700496 348851 700498
rect 292481 700440 292486 700496
rect 292542 700440 348790 700496
rect 348846 700440 348851 700496
rect 292481 700438 348851 700440
rect 292481 700435 292547 700438
rect 348785 700435 348851 700438
rect 296478 700300 296484 700364
rect 296548 700362 296554 700364
rect 413645 700362 413711 700365
rect 296548 700360 413711 700362
rect 296548 700304 413650 700360
rect 413706 700304 413711 700360
rect 296548 700302 413711 700304
rect 296548 700300 296554 700302
rect 413645 700299 413711 700302
rect 559649 700362 559715 700365
rect 582373 700362 582439 700365
rect 559649 700360 582439 700362
rect 559649 700304 559654 700360
rect 559710 700304 582378 700360
rect 582434 700304 582439 700360
rect 559649 700302 582439 700304
rect 559649 700299 559715 700302
rect 582373 700299 582439 700302
rect 289721 697506 289787 697509
rect 478505 697506 478571 697509
rect 289721 697504 478571 697506
rect -960 697220 480 697460
rect 289721 697448 289726 697504
rect 289782 697448 478510 697504
rect 478566 697448 478571 697504
rect 289721 697446 478571 697448
rect 289721 697443 289787 697446
rect 478505 697443 478571 697446
rect 543457 697506 543523 697509
rect 543457 697504 567210 697506
rect 543457 697448 543462 697504
rect 543518 697448 567210 697504
rect 543457 697446 567210 697448
rect 543457 697443 543523 697446
rect 567150 697234 567210 697446
rect 580901 697234 580967 697237
rect 583520 697234 584960 697324
rect 567150 697232 584960 697234
rect 567150 697176 580906 697232
rect 580962 697176 584960 697232
rect 567150 697174 584960 697176
rect 580901 697171 580967 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 8886 684314 8892 684316
rect -960 684254 8892 684314
rect -960 684164 480 684254
rect 8886 684252 8892 684254
rect 8956 684252 8962 684316
rect 580901 683906 580967 683909
rect 583520 683906 584960 683996
rect 580901 683904 584960 683906
rect 580901 683848 580906 683904
rect 580962 683848 584960 683904
rect 580901 683846 584960 683848
rect 580901 683843 580967 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 285622 671258 285628 671260
rect -960 671198 285628 671258
rect -960 671108 480 671198
rect 285622 671196 285628 671198
rect 285692 671196 285698 671260
rect 575974 670652 575980 670716
rect 576044 670714 576050 670716
rect 583520 670714 584960 670804
rect 576044 670654 584960 670714
rect 576044 670652 576050 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 290406 658202 290412 658204
rect -960 658142 290412 658202
rect -960 658052 480 658142
rect 290406 658140 290412 658142
rect 290476 658140 290482 658204
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580901 644058 580967 644061
rect 583520 644058 584960 644148
rect 580901 644056 584960 644058
rect 580901 644000 580906 644056
rect 580962 644000 584960 644056
rect 580901 643998 584960 644000
rect 580901 643995 580967 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 1894 632090 1900 632092
rect -960 632030 1900 632090
rect -960 631940 480 632030
rect 1894 632028 1900 632030
rect 1964 632028 1970 632092
rect 580901 630866 580967 630869
rect 583520 630866 584960 630956
rect 580901 630864 584960 630866
rect 580901 630808 580906 630864
rect 580962 630808 584960 630864
rect 580901 630806 584960 630808
rect 580901 630803 580967 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 281022 619170 281028 619172
rect -960 619110 281028 619170
rect -960 619020 480 619110
rect 281022 619108 281028 619110
rect 281092 619108 281098 619172
rect 576158 617476 576164 617540
rect 576228 617538 576234 617540
rect 583520 617538 584960 617628
rect 576228 617478 584960 617538
rect 576228 617476 576234 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect -960 606054 674 606114
rect -960 605978 480 606054
rect 614 605978 674 606054
rect -960 605964 674 605978
rect 62 605918 674 605964
rect 62 605844 122 605918
rect 54 605780 60 605844
rect 124 605780 130 605844
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580901 591018 580967 591021
rect 583520 591018 584960 591108
rect 580901 591016 584960 591018
rect 580901 590960 580906 591016
rect 580962 590960 584960 591016
rect 580901 590958 584960 590960
rect 580901 590955 580967 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 4654 580002 4660 580004
rect -960 579942 4660 580002
rect -960 579852 480 579942
rect 4654 579940 4660 579942
rect 4724 579940 4730 580004
rect 580901 577690 580967 577693
rect 583520 577690 584960 577780
rect 580901 577688 584960 577690
rect 580901 577632 580906 577688
rect 580962 577632 584960 577688
rect 580901 577630 584960 577632
rect 580901 577627 580967 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 7414 566946 7420 566948
rect -960 566886 7420 566946
rect -960 566796 480 566886
rect 7414 566884 7420 566886
rect 7484 566884 7490 566948
rect 574686 564300 574692 564364
rect 574756 564362 574762 564364
rect 583520 564362 584960 564452
rect 574756 564302 584960 564362
rect 574756 564300 574762 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 4838 553890 4844 553892
rect -960 553830 4844 553890
rect -960 553740 480 553830
rect 4838 553828 4844 553830
rect 4908 553828 4914 553892
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580901 537842 580967 537845
rect 583520 537842 584960 537932
rect 580901 537840 584960 537842
rect 580901 537784 580906 537840
rect 580962 537784 584960 537840
rect 580901 537782 584960 537784
rect 580901 537779 580967 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 9070 527914 9076 527916
rect -960 527854 9076 527914
rect -960 527764 480 527854
rect 9070 527852 9076 527854
rect 9140 527852 9146 527916
rect 580901 524514 580967 524517
rect 583520 524514 584960 524604
rect 580901 524512 584960 524514
rect 580901 524456 580906 524512
rect 580962 524456 584960 524512
rect 580901 524454 584960 524456
rect 580901 524451 580967 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 6126 514858 6132 514860
rect -960 514798 6132 514858
rect -960 514708 480 514798
rect 6126 514796 6132 514798
rect 6196 514796 6202 514860
rect 574870 511260 574876 511324
rect 574940 511322 574946 511324
rect 583520 511322 584960 511412
rect 574940 511262 584960 511322
rect 574940 511260 574946 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 7598 501802 7604 501804
rect -960 501742 7604 501802
rect -960 501652 480 501742
rect 7598 501740 7604 501742
rect 7668 501740 7674 501804
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580901 484666 580967 484669
rect 583520 484666 584960 484756
rect 580901 484664 584960 484666
rect 580901 484608 580906 484664
rect 580962 484608 584960 484664
rect 580901 484606 584960 484608
rect 580901 484603 580967 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 7782 475690 7788 475692
rect -960 475630 7788 475690
rect -960 475540 480 475630
rect 7782 475628 7788 475630
rect 7852 475628 7858 475692
rect 580901 471474 580967 471477
rect 583520 471474 584960 471564
rect 580901 471472 584960 471474
rect 580901 471416 580906 471472
rect 580962 471416 584960 471472
rect 580901 471414 584960 471416
rect 580901 471411 580967 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 12382 462634 12388 462636
rect -960 462574 12388 462634
rect -960 462484 480 462574
rect 12382 462572 12388 462574
rect 12452 462572 12458 462636
rect 578734 458084 578740 458148
rect 578804 458146 578810 458148
rect 583520 458146 584960 458236
rect 578804 458086 584960 458146
rect 578804 458084 578810 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 6310 449578 6316 449580
rect -960 449518 6316 449578
rect -960 449428 480 449518
rect 6310 449516 6316 449518
rect 6380 449516 6386 449580
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580901 431626 580967 431629
rect 583520 431626 584960 431716
rect 580901 431624 584960 431626
rect 580901 431568 580906 431624
rect 580962 431568 584960 431624
rect 580901 431566 584960 431568
rect 580901 431563 580967 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 9254 423602 9260 423604
rect -960 423542 9260 423602
rect -960 423452 480 423542
rect 9254 423540 9260 423542
rect 9324 423540 9330 423604
rect 580901 418298 580967 418301
rect 583520 418298 584960 418388
rect 580901 418296 584960 418298
rect 580901 418240 580906 418296
rect 580962 418240 584960 418296
rect 580901 418238 584960 418240
rect 580901 418235 580967 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 11094 410546 11100 410548
rect -960 410486 11100 410546
rect -960 410396 480 410486
rect 11094 410484 11100 410486
rect 11164 410484 11170 410548
rect 577446 404908 577452 404972
rect 577516 404970 577522 404972
rect 583520 404970 584960 405060
rect 577516 404910 584960 404970
rect 577516 404908 577522 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 6494 397490 6500 397492
rect -960 397430 6500 397490
rect -960 397340 480 397430
rect 6494 397428 6500 397430
rect 6564 397428 6570 397492
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580901 378450 580967 378453
rect 583520 378450 584960 378540
rect 580901 378448 584960 378450
rect 580901 378392 580906 378448
rect 580962 378392 584960 378448
rect 580901 378390 584960 378392
rect 580901 378387 580967 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 9806 371378 9812 371380
rect -960 371318 9812 371378
rect -960 371228 480 371318
rect 9806 371316 9812 371318
rect 9876 371316 9882 371380
rect 580901 365122 580967 365125
rect 583520 365122 584960 365212
rect 580901 365120 584960 365122
rect 580901 365064 580906 365120
rect 580962 365064 584960 365120
rect 580901 365062 584960 365064
rect 580901 365059 580967 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3366 358458 3372 358460
rect -960 358398 3372 358458
rect -960 358308 480 358398
rect 3366 358396 3372 358398
rect 3436 358396 3442 358460
rect 577630 351868 577636 351932
rect 577700 351930 577706 351932
rect 583520 351930 584960 352020
rect 577700 351870 584960 351930
rect 577700 351868 577706 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 2078 345402 2084 345404
rect -960 345342 2084 345402
rect -960 345252 480 345342
rect 2078 345340 2084 345342
rect 2148 345340 2154 345404
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580901 325274 580967 325277
rect 583520 325274 584960 325364
rect 580901 325272 584960 325274
rect 580901 325216 580906 325272
rect 580962 325216 584960 325272
rect 580901 325214 584960 325216
rect 580901 325211 580967 325214
rect 583520 325124 584960 325214
rect 420952 323444 420958 323508
rect 421022 323506 421028 323508
rect 422176 323506 422182 323508
rect 421022 323446 422182 323506
rect 421022 323444 421028 323446
rect 422176 323444 422182 323446
rect 422246 323506 422252 323508
rect 433328 323506 433334 323508
rect 422246 323444 422310 323506
rect 422250 323370 422310 323444
rect 431910 323446 433334 323506
rect 431910 323370 431970 323446
rect 433328 323444 433334 323446
rect 433398 323506 433404 323508
rect 439129 323506 439195 323509
rect 433398 323504 439195 323506
rect 433398 323448 439134 323504
rect 439190 323448 439195 323504
rect 433398 323446 439195 323448
rect 433398 323444 433404 323446
rect 439129 323443 439195 323446
rect 422250 323310 431970 323370
rect 439129 319834 439195 319837
rect 439086 319832 439195 319834
rect 439086 319776 439134 319832
rect 439190 319776 439195 319832
rect 439086 319771 439195 319776
rect 439086 319426 439146 319771
rect -960 319290 480 319380
rect 439086 319366 439514 319426
rect 3550 319290 3556 319292
rect -960 319230 3556 319290
rect -960 319140 480 319230
rect 3550 319228 3556 319230
rect 3620 319228 3626 319292
rect 439454 319290 439514 319366
rect 441654 319290 441660 319292
rect 439454 319230 441660 319290
rect 439454 319220 439514 319230
rect 441654 319228 441660 319230
rect 441724 319228 441730 319292
rect 439116 319160 439514 319220
rect 580901 312082 580967 312085
rect 583520 312082 584960 312172
rect 580901 312080 584960 312082
rect 580901 312024 580906 312080
rect 580962 312024 584960 312080
rect 580901 312022 584960 312024
rect 580901 312019 580967 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3734 306234 3740 306236
rect -960 306174 3740 306234
rect -960 306084 480 306174
rect 3734 306172 3740 306174
rect 3804 306172 3810 306236
rect 580206 298692 580212 298756
rect 580276 298754 580282 298756
rect 583520 298754 584960 298844
rect 580276 298694 584960 298754
rect 580276 298692 580282 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect -960 293118 674 293178
rect -960 293042 480 293118
rect 614 293042 674 293118
rect -960 293028 674 293042
rect 246 292982 674 293028
rect 246 292636 306 292982
rect 238 292572 244 292636
rect 308 292572 314 292636
rect 583520 285276 584960 285516
rect 154113 281074 154179 281077
rect 281942 281074 281948 281076
rect 154113 281072 281948 281074
rect 154113 281016 154118 281072
rect 154174 281016 281948 281072
rect 154113 281014 281948 281016
rect 154113 281011 154179 281014
rect 281942 281012 281948 281014
rect 282012 281012 282018 281076
rect 89161 280938 89227 280941
rect 287094 280938 287100 280940
rect 89161 280936 287100 280938
rect 89161 280880 89166 280936
rect 89222 280880 287100 280936
rect 89161 280878 287100 280880
rect 89161 280875 89227 280878
rect 287094 280876 287100 280878
rect 287164 280876 287170 280940
rect 24301 280802 24367 280805
rect 284334 280802 284340 280804
rect 24301 280800 284340 280802
rect 24301 280744 24306 280800
rect 24362 280744 284340 280800
rect 24301 280742 284340 280744
rect 24301 280739 24367 280742
rect 284334 280740 284340 280742
rect 284404 280740 284410 280804
rect -960 279972 480 280212
rect 301822 276864 302496 276924
rect 300526 276796 300532 276860
rect 300596 276858 300602 276860
rect 301822 276858 301882 276864
rect 300596 276798 301882 276858
rect 300596 276796 300602 276798
rect 301998 275910 302004 275974
rect 302068 275972 302074 275974
rect 302068 275912 302496 275972
rect 302068 275910 302074 275912
rect 302006 273736 302496 273796
rect 301814 273668 301820 273732
rect 301884 273730 301890 273732
rect 302006 273730 302066 273736
rect 301884 273670 302066 273730
rect 301884 273668 301890 273670
rect 301822 272784 302496 272844
rect 301630 272716 301636 272780
rect 301700 272778 301706 272780
rect 301822 272778 301882 272784
rect 301700 272718 301882 272778
rect 301700 272716 301706 272718
rect 580901 272234 580967 272237
rect 583520 272234 584960 272324
rect 580901 272232 584960 272234
rect 580901 272176 580906 272232
rect 580962 272176 584960 272232
rect 580901 272174 584960 272176
rect 580901 272171 580967 272174
rect 583520 272084 584960 272174
rect 3550 271764 3556 271828
rect 3620 271826 3626 271828
rect 5022 271826 5028 271828
rect 3620 271766 5028 271826
rect 3620 271764 3626 271766
rect 5022 271764 5028 271766
rect 5092 271764 5098 271828
rect 301822 271016 302496 271076
rect 300710 270948 300716 271012
rect 300780 271010 300786 271012
rect 301822 271010 301882 271016
rect 300780 270950 301882 271010
rect 300780 270948 300786 270950
rect 301822 269928 302496 269988
rect 300158 269860 300164 269924
rect 300228 269922 300234 269924
rect 301822 269922 301882 269928
rect 300228 269862 301882 269922
rect 300228 269860 300234 269862
rect 301822 268160 302496 268220
rect 300342 268092 300348 268156
rect 300412 268154 300418 268156
rect 301822 268154 301882 268160
rect 300412 268094 301882 268154
rect 300412 268092 300418 268094
rect -960 267202 480 267292
rect 3550 267202 3556 267204
rect -960 267142 3556 267202
rect -960 267052 480 267142
rect 3550 267140 3556 267142
rect 3620 267140 3626 267204
rect 439270 259390 439698 259450
rect 439270 259380 439330 259390
rect 439116 259320 439330 259380
rect 439638 259314 439698 259390
rect 580574 259388 580580 259452
rect 580644 259450 580650 259452
rect 580901 259450 580967 259453
rect 580644 259448 580967 259450
rect 580644 259392 580906 259448
rect 580962 259392 580967 259448
rect 580644 259390 580967 259392
rect 580644 259388 580650 259390
rect 580901 259387 580967 259390
rect 441654 259314 441660 259316
rect 439638 259254 441660 259314
rect 439638 259178 439698 259254
rect 441654 259252 441660 259254
rect 441724 259252 441730 259316
rect 439086 259118 439698 259178
rect 439086 257954 439146 259118
rect 580574 258844 580580 258908
rect 580644 258906 580650 258908
rect 583520 258906 584960 258996
rect 580644 258846 584960 258906
rect 580644 258844 580650 258846
rect 583520 258756 584960 258846
rect 439086 257894 439514 257954
rect 439454 257748 439514 257894
rect 439116 257688 439514 257748
rect 439454 257546 439514 257688
rect 439086 257486 439514 257546
rect 439086 256594 439146 257486
rect 439086 256534 439514 256594
rect 439454 256388 439514 256534
rect 439116 256328 439514 256388
rect 439454 256186 439514 256328
rect 439086 256126 439514 256186
rect 439086 255098 439146 256126
rect 439086 255038 439514 255098
rect 439454 254892 439514 255038
rect 439116 254832 439514 254892
rect 439454 254690 439514 254832
rect 439086 254630 439514 254690
rect -960 254146 480 254236
rect -960 254086 2146 254146
rect -960 253996 480 254086
rect 2086 254010 2146 254086
rect 2773 254010 2839 254013
rect 3417 254010 3483 254013
rect 2086 254008 3483 254010
rect 2086 253952 2778 254008
rect 2834 253952 3422 254008
rect 3478 253952 3483 254008
rect 2086 253950 3483 253952
rect 2773 253947 2839 253950
rect 3417 253947 3483 253950
rect 439086 253874 439146 254630
rect 439086 253814 439514 253874
rect 439116 253608 439330 253668
rect 439270 253602 439330 253608
rect 439454 253602 439514 253814
rect 441654 253602 441660 253604
rect 439270 253542 441660 253602
rect 441654 253540 441660 253542
rect 441724 253540 441730 253604
rect 301822 249936 302496 249996
rect 301446 249868 301452 249932
rect 301516 249930 301522 249932
rect 301822 249930 301882 249936
rect 301516 249870 301882 249930
rect 301516 249868 301522 249870
rect 300526 249732 300532 249796
rect 300596 249794 300602 249796
rect 302366 249794 302372 249796
rect 300596 249734 302372 249794
rect 300596 249732 300602 249734
rect 302366 249732 302372 249734
rect 302436 249732 302442 249796
rect 301822 248304 302496 248364
rect 299974 248236 299980 248300
rect 300044 248298 300050 248300
rect 301822 248298 301882 248304
rect 300044 248238 301882 248298
rect 300044 248236 300050 248238
rect 301822 248032 302496 248092
rect 300526 247964 300532 248028
rect 300596 248026 300602 248028
rect 301822 248026 301882 248032
rect 300596 247966 301882 248026
rect 300596 247964 300602 247966
rect 300158 247012 300164 247076
rect 300228 247074 300234 247076
rect 300761 247074 300827 247077
rect 300228 247072 300827 247074
rect 300228 247016 300766 247072
rect 300822 247016 300827 247072
rect 300228 247014 300827 247016
rect 300228 247012 300234 247014
rect 300761 247011 300827 247014
rect 578918 245516 578924 245580
rect 578988 245578 578994 245580
rect 583520 245578 584960 245668
rect 578988 245518 584960 245578
rect 578988 245516 578994 245518
rect 583520 245428 584960 245518
rect 3734 242796 3740 242860
rect 3804 242858 3810 242860
rect 9438 242858 9444 242860
rect 3804 242798 9444 242858
rect 3804 242796 3810 242798
rect 9438 242796 9444 242798
rect 9508 242796 9514 242860
rect -960 241090 480 241180
rect 2814 241090 2820 241092
rect -960 241030 2820 241090
rect -960 240940 480 241030
rect 2814 241028 2820 241030
rect 2884 241028 2890 241092
rect 301446 239940 301452 240004
rect 301516 240002 301522 240004
rect 304758 240002 304764 240004
rect 301516 239942 304764 240002
rect 301516 239940 301522 239942
rect 304758 239940 304764 239942
rect 304828 239940 304834 240004
rect 441654 240002 441660 240004
rect 425856 239942 441660 240002
rect 425856 239868 425916 239942
rect 441654 239940 441660 239942
rect 441724 239940 441730 240004
rect 425848 239804 425854 239868
rect 425918 239804 425924 239868
rect 337326 237900 337332 237964
rect 337396 237962 337402 237964
rect 425830 237962 425836 237964
rect 337396 237902 425836 237962
rect 337396 237900 337402 237902
rect 425830 237900 425836 237902
rect 425900 237900 425906 237964
rect 300342 237356 300348 237420
rect 300412 237418 300418 237420
rect 308254 237418 308260 237420
rect 300412 237358 308260 237418
rect 300412 237356 300418 237358
rect 308254 237356 308260 237358
rect 308324 237356 308330 237420
rect 329414 236812 329420 236876
rect 329484 236874 329490 236876
rect 353334 236874 353340 236876
rect 329484 236814 353340 236874
rect 329484 236812 329490 236814
rect 353334 236812 353340 236814
rect 353404 236812 353410 236876
rect 312486 236676 312492 236740
rect 312556 236738 312562 236740
rect 324262 236738 324268 236740
rect 312556 236678 324268 236738
rect 312556 236676 312562 236678
rect 324262 236676 324268 236678
rect 324332 236676 324338 236740
rect 325366 236676 325372 236740
rect 325436 236738 325442 236740
rect 350758 236738 350764 236740
rect 325436 236678 350764 236738
rect 325436 236676 325442 236678
rect 350758 236676 350764 236678
rect 350828 236676 350834 236740
rect 323526 236540 323532 236604
rect 323596 236602 323602 236604
rect 336958 236602 336964 236604
rect 323596 236542 336964 236602
rect 323596 236540 323602 236542
rect 336958 236540 336964 236542
rect 337028 236540 337034 236604
rect 349654 236540 349660 236604
rect 349724 236602 349730 236604
rect 408350 236602 408356 236604
rect 349724 236542 408356 236602
rect 349724 236540 349730 236542
rect 408350 236540 408356 236542
rect 408420 236540 408426 236604
rect 337878 236132 337884 236196
rect 337948 236194 337954 236196
rect 340454 236194 340460 236196
rect 337948 236134 340460 236194
rect 337948 236132 337954 236134
rect 340454 236132 340460 236134
rect 340524 236132 340530 236196
rect 299974 235996 299980 236060
rect 300044 236058 300050 236060
rect 305678 236058 305684 236060
rect 300044 235998 305684 236058
rect 300044 235996 300050 235998
rect 305678 235996 305684 235998
rect 305748 235996 305754 236060
rect 316534 235996 316540 236060
rect 316604 236058 316610 236060
rect 318558 236058 318564 236060
rect 316604 235998 318564 236058
rect 316604 235996 316610 235998
rect 318558 235996 318564 235998
rect 318628 235996 318634 236060
rect 319478 235996 319484 236060
rect 319548 236058 319554 236060
rect 322974 236058 322980 236060
rect 319548 235998 322980 236058
rect 319548 235996 319554 235998
rect 322974 235996 322980 235998
rect 323044 235996 323050 236060
rect 323158 235996 323164 236060
rect 323228 236058 323234 236060
rect 325550 236058 325556 236060
rect 323228 235998 325556 236058
rect 323228 235996 323234 235998
rect 325550 235996 325556 235998
rect 325620 235996 325626 236060
rect 334566 235996 334572 236060
rect 334636 236058 334642 236060
rect 336222 236058 336228 236060
rect 334636 235998 336228 236058
rect 334636 235996 334642 235998
rect 336222 235996 336228 235998
rect 336292 235996 336298 236060
rect 340270 235996 340276 236060
rect 340340 236058 340346 236060
rect 344134 236058 344140 236060
rect 340340 235998 344140 236058
rect 340340 235996 340346 235998
rect 344134 235996 344140 235998
rect 344204 235996 344210 236060
rect 300710 235860 300716 235924
rect 300780 235922 300786 235924
rect 308990 235922 308996 235924
rect 300780 235862 308996 235922
rect 300780 235860 300786 235862
rect 308990 235860 308996 235862
rect 309060 235860 309066 235924
rect 323710 235588 323716 235652
rect 323780 235650 323786 235652
rect 338614 235650 338620 235652
rect 323780 235590 338620 235650
rect 323780 235588 323786 235590
rect 338614 235588 338620 235590
rect 338684 235588 338690 235652
rect 313406 235452 313412 235516
rect 313476 235514 313482 235516
rect 333830 235514 333836 235516
rect 313476 235454 333836 235514
rect 313476 235452 313482 235454
rect 333830 235452 333836 235454
rect 333900 235452 333906 235516
rect 333094 235316 333100 235380
rect 333164 235378 333170 235380
rect 366030 235378 366036 235380
rect 333164 235318 366036 235378
rect 333164 235316 333170 235318
rect 366030 235316 366036 235318
rect 366100 235316 366106 235380
rect 320766 235180 320772 235244
rect 320836 235242 320842 235244
rect 356830 235242 356836 235244
rect 320836 235182 356836 235242
rect 320836 235180 320842 235182
rect 356830 235180 356836 235182
rect 356900 235180 356906 235244
rect 324998 234092 325004 234156
rect 325068 234154 325074 234156
rect 343214 234154 343220 234156
rect 325068 234094 343220 234154
rect 325068 234092 325074 234094
rect 343214 234092 343220 234094
rect 343284 234092 343290 234156
rect 78438 233956 78444 234020
rect 78508 234018 78514 234020
rect 90030 234018 90036 234020
rect 78508 233958 90036 234018
rect 78508 233956 78514 233958
rect 90030 233956 90036 233958
rect 90100 233956 90106 234020
rect 318558 233956 318564 234020
rect 318628 234018 318634 234020
rect 350022 234018 350028 234020
rect 318628 233958 350028 234018
rect 318628 233956 318634 233958
rect 350022 233956 350028 233958
rect 350092 233956 350098 234020
rect 89294 233820 89300 233884
rect 89364 233882 89370 233884
rect 110454 233882 110460 233884
rect 89364 233822 110460 233882
rect 89364 233820 89370 233822
rect 110454 233820 110460 233822
rect 110524 233820 110530 233884
rect 301630 233820 301636 233884
rect 301700 233882 301706 233884
rect 309358 233882 309364 233884
rect 301700 233822 309364 233882
rect 301700 233820 301706 233822
rect 309358 233820 309364 233822
rect 309428 233820 309434 233884
rect 310830 233820 310836 233884
rect 310900 233882 310906 233884
rect 323158 233882 323164 233884
rect 310900 233822 323164 233882
rect 310900 233820 310906 233822
rect 323158 233820 323164 233822
rect 323228 233820 323234 233884
rect 327390 233820 327396 233884
rect 327460 233882 327466 233884
rect 363454 233882 363460 233884
rect 327460 233822 363460 233882
rect 327460 233820 327466 233822
rect 363454 233820 363460 233822
rect 363524 233820 363530 233884
rect 317454 232732 317460 232796
rect 317524 232794 317530 232796
rect 346342 232794 346348 232796
rect 317524 232734 346348 232794
rect 317524 232732 317530 232734
rect 346342 232732 346348 232734
rect 346412 232732 346418 232796
rect 321870 232596 321876 232660
rect 321940 232658 321946 232660
rect 360510 232658 360516 232660
rect 321940 232598 360516 232658
rect 321940 232596 321946 232598
rect 360510 232596 360516 232598
rect 360580 232596 360586 232660
rect 301814 232460 301820 232524
rect 301884 232522 301890 232524
rect 309726 232522 309732 232524
rect 301884 232462 309732 232522
rect 301884 232460 301890 232462
rect 309726 232460 309732 232462
rect 309796 232460 309802 232524
rect 314878 232460 314884 232524
rect 314948 232522 314954 232524
rect 338246 232522 338252 232524
rect 314948 232462 338252 232522
rect 314948 232460 314954 232462
rect 338246 232460 338252 232462
rect 338316 232460 338322 232524
rect 338614 232460 338620 232524
rect 338684 232522 338690 232524
rect 400990 232522 400996 232524
rect 338684 232462 400996 232522
rect 338684 232460 338690 232462
rect 400990 232460 400996 232462
rect 401060 232460 401066 232524
rect 580901 232386 580967 232389
rect 583520 232386 584960 232476
rect 580901 232384 584960 232386
rect 580901 232328 580906 232384
rect 580962 232328 584960 232384
rect 580901 232326 584960 232328
rect 580901 232323 580967 232326
rect 583520 232236 584960 232326
rect 315614 231372 315620 231436
rect 315684 231434 315690 231436
rect 337878 231434 337884 231436
rect 315684 231374 337884 231434
rect 315684 231372 315690 231374
rect 337878 231372 337884 231374
rect 337948 231372 337954 231436
rect 318190 231236 318196 231300
rect 318260 231298 318266 231300
rect 348918 231298 348924 231300
rect 318260 231238 348924 231298
rect 318260 231236 318266 231238
rect 348918 231236 348924 231238
rect 348988 231236 348994 231300
rect 360694 231236 360700 231300
rect 360764 231298 360770 231300
rect 370814 231298 370820 231300
rect 360764 231238 370820 231298
rect 360764 231236 360770 231238
rect 370814 231236 370820 231238
rect 370884 231236 370890 231300
rect 326654 231100 326660 231164
rect 326724 231162 326730 231164
rect 361062 231162 361068 231164
rect 326724 231102 361068 231162
rect 326724 231100 326730 231102
rect 361062 231100 361068 231102
rect 361132 231100 361138 231164
rect 326470 230420 326476 230484
rect 326540 230482 326546 230484
rect 333278 230482 333284 230484
rect 326540 230422 333284 230482
rect 326540 230420 326546 230422
rect 333278 230420 333284 230422
rect 333348 230420 333354 230484
rect 315798 230012 315804 230076
rect 315868 230074 315874 230076
rect 342110 230074 342116 230076
rect 315868 230014 342116 230074
rect 315868 230012 315874 230014
rect 342110 230012 342116 230014
rect 342180 230012 342186 230076
rect 321134 229876 321140 229940
rect 321204 229938 321210 229940
rect 358302 229938 358308 229940
rect 321204 229878 358308 229938
rect 321204 229876 321210 229878
rect 358302 229876 358308 229878
rect 358372 229876 358378 229940
rect 306046 229740 306052 229804
rect 306116 229802 306122 229804
rect 320582 229802 320588 229804
rect 306116 229742 320588 229802
rect 306116 229740 306122 229742
rect 320582 229740 320588 229742
rect 320652 229740 320658 229804
rect 333646 229740 333652 229804
rect 333716 229802 333722 229804
rect 405590 229802 405596 229804
rect 333716 229742 405596 229802
rect 333716 229740 333722 229742
rect 405590 229740 405596 229742
rect 405660 229740 405666 229804
rect 315246 228516 315252 228580
rect 315316 228578 315322 228580
rect 339534 228578 339540 228580
rect 315316 228518 339540 228578
rect 315316 228516 315322 228518
rect 339534 228516 339540 228518
rect 339604 228516 339610 228580
rect 327574 228380 327580 228444
rect 327644 228442 327650 228444
rect 356094 228442 356100 228444
rect 327644 228382 356100 228442
rect 327644 228380 327650 228382
rect 356094 228380 356100 228382
rect 356164 228380 356170 228444
rect 317822 228244 317828 228308
rect 317892 228306 317898 228308
rect 347814 228306 347820 228308
rect 317892 228246 347820 228306
rect 317892 228244 317898 228246
rect 347814 228244 347820 228246
rect 347884 228244 347890 228308
rect 356646 228244 356652 228308
rect 356716 228306 356722 228308
rect 395838 228306 395844 228308
rect 356716 228246 395844 228306
rect 356716 228244 356722 228246
rect 395838 228244 395844 228246
rect 395908 228244 395914 228308
rect -960 227884 480 228124
rect 317086 227156 317092 227220
rect 317156 227218 317162 227220
rect 345422 227218 345428 227220
rect 317156 227158 345428 227218
rect 317156 227156 317162 227158
rect 345422 227156 345428 227158
rect 345492 227156 345498 227220
rect 321318 227020 321324 227084
rect 321388 227082 321394 227084
rect 359590 227082 359596 227084
rect 321388 227022 359596 227082
rect 321388 227020 321394 227022
rect 359590 227020 359596 227022
rect 359660 227020 359666 227084
rect 314510 226884 314516 226948
rect 314580 226946 314586 226948
rect 323526 226946 323532 226948
rect 314580 226886 323532 226946
rect 314580 226884 314586 226886
rect 323526 226884 323532 226886
rect 323596 226884 323602 226948
rect 331990 226884 331996 226948
rect 332060 226946 332066 226948
rect 386086 226946 386092 226948
rect 332060 226886 386092 226946
rect 332060 226884 332066 226886
rect 386086 226884 386092 226886
rect 386156 226884 386162 226948
rect 311934 225932 311940 225996
rect 312004 225994 312010 225996
rect 329046 225994 329052 225996
rect 312004 225934 329052 225994
rect 312004 225932 312010 225934
rect 329046 225932 329052 225934
rect 329116 225932 329122 225996
rect 340086 225932 340092 225996
rect 340156 225994 340162 225996
rect 348550 225994 348556 225996
rect 340156 225934 348556 225994
rect 340156 225932 340162 225934
rect 348550 225932 348556 225934
rect 348620 225932 348626 225996
rect 324814 225796 324820 225860
rect 324884 225858 324890 225860
rect 346158 225858 346164 225860
rect 324884 225798 346164 225858
rect 324884 225796 324890 225798
rect 346158 225796 346164 225798
rect 346228 225796 346234 225860
rect 316718 225660 316724 225724
rect 316788 225722 316794 225724
rect 340270 225722 340276 225724
rect 316788 225662 340276 225722
rect 316788 225660 316794 225662
rect 340270 225660 340276 225662
rect 340340 225660 340346 225724
rect 328494 225524 328500 225588
rect 328564 225586 328570 225588
rect 368606 225586 368612 225588
rect 328564 225526 368612 225586
rect 328564 225524 328570 225526
rect 368606 225524 368612 225526
rect 368676 225524 368682 225588
rect 307150 224980 307156 225044
rect 307220 225042 307226 225044
rect 312486 225042 312492 225044
rect 307220 224982 312492 225042
rect 307220 224980 307226 224982
rect 312486 224980 312492 224982
rect 312556 224980 312562 225044
rect 324078 224436 324084 224500
rect 324148 224498 324154 224500
rect 341006 224498 341012 224500
rect 324148 224438 341012 224498
rect 324148 224436 324154 224438
rect 341006 224436 341012 224438
rect 341076 224436 341082 224500
rect 307886 224300 307892 224364
rect 307956 224362 307962 224364
rect 319662 224362 319668 224364
rect 307956 224302 319668 224362
rect 307956 224300 307962 224302
rect 319662 224300 319668 224302
rect 319732 224300 319738 224364
rect 331438 224300 331444 224364
rect 331508 224362 331514 224364
rect 391054 224362 391060 224364
rect 331508 224302 391060 224362
rect 331508 224300 331514 224302
rect 391054 224300 391060 224302
rect 391124 224300 391130 224364
rect 312486 224164 312492 224228
rect 312556 224226 312562 224228
rect 327942 224226 327948 224228
rect 312556 224166 327948 224226
rect 312556 224164 312562 224166
rect 327942 224164 327948 224166
rect 328012 224164 328018 224228
rect 328310 224164 328316 224228
rect 328380 224226 328386 224228
rect 331254 224226 331260 224228
rect 328380 224166 331260 224226
rect 328380 224164 328386 224166
rect 331254 224164 331260 224166
rect 331324 224164 331330 224228
rect 332358 224164 332364 224228
rect 332428 224226 332434 224228
rect 398414 224226 398420 224228
rect 332428 224166 398420 224226
rect 332428 224164 332434 224166
rect 398414 224164 398420 224166
rect 398484 224164 398490 224228
rect 322606 223212 322612 223276
rect 322676 223274 322682 223276
rect 330886 223274 330892 223276
rect 322676 223214 330892 223274
rect 322676 223212 322682 223214
rect 330886 223212 330892 223214
rect 330956 223212 330962 223276
rect 330518 223076 330524 223140
rect 330588 223138 330594 223140
rect 343582 223138 343588 223140
rect 330588 223078 343588 223138
rect 330588 223076 330594 223078
rect 343582 223076 343588 223078
rect 343652 223076 343658 223140
rect 323342 222940 323348 223004
rect 323412 223002 323418 223004
rect 334566 223002 334572 223004
rect 323412 222942 334572 223002
rect 323412 222940 323418 222942
rect 334566 222940 334572 222942
rect 334636 222940 334642 223004
rect 334750 222940 334756 223004
rect 334820 223002 334826 223004
rect 373574 223002 373580 223004
rect 334820 222942 373580 223002
rect 334820 222940 334826 222942
rect 373574 222940 373580 222942
rect 373644 222940 373650 223004
rect 311014 222804 311020 222868
rect 311084 222866 311090 222868
rect 322238 222866 322244 222868
rect 311084 222806 322244 222866
rect 311084 222804 311090 222806
rect 322238 222804 322244 222806
rect 322308 222804 322314 222868
rect 330334 222804 330340 222868
rect 330404 222866 330410 222868
rect 383510 222866 383516 222868
rect 330404 222806 383516 222866
rect 330404 222804 330410 222806
rect 383510 222804 383516 222806
rect 383580 222804 383586 222868
rect 334566 221852 334572 221916
rect 334636 221914 334642 221916
rect 349654 221914 349660 221916
rect 334636 221854 349660 221914
rect 334636 221852 334642 221854
rect 349654 221852 349660 221854
rect 349724 221852 349730 221916
rect 313774 221716 313780 221780
rect 313844 221778 313850 221780
rect 334934 221778 334940 221780
rect 313844 221718 334940 221778
rect 313844 221716 313850 221718
rect 334934 221716 334940 221718
rect 335004 221716 335010 221780
rect 322238 221580 322244 221644
rect 322308 221642 322314 221644
rect 361798 221642 361804 221644
rect 322308 221582 361804 221642
rect 322308 221580 322314 221582
rect 361798 221580 361804 221582
rect 361868 221580 361874 221644
rect 313038 221444 313044 221508
rect 313108 221506 313114 221508
rect 332726 221506 332732 221508
rect 313108 221446 332732 221506
rect 313108 221444 313114 221446
rect 332726 221444 332732 221446
rect 332796 221444 332802 221508
rect 333278 221444 333284 221508
rect 333348 221506 333354 221508
rect 403566 221506 403572 221508
rect 333348 221446 403572 221506
rect 333348 221444 333354 221446
rect 403566 221444 403572 221446
rect 403636 221444 403642 221508
rect 300761 220962 300827 220965
rect 307753 220962 307819 220965
rect 300761 220960 307819 220962
rect 300761 220904 300766 220960
rect 300822 220904 307758 220960
rect 307814 220904 307819 220960
rect 300761 220902 307819 220904
rect 300761 220899 300827 220902
rect 307753 220899 307819 220902
rect 320030 220356 320036 220420
rect 320100 220418 320106 220420
rect 354438 220418 354444 220420
rect 320100 220358 354444 220418
rect 320100 220356 320106 220358
rect 354438 220356 354444 220358
rect 354508 220356 354514 220420
rect 320398 220220 320404 220284
rect 320468 220282 320474 220284
rect 355910 220282 355916 220284
rect 320468 220222 355916 220282
rect 320468 220220 320474 220222
rect 355910 220220 355916 220222
rect 355980 220220 355986 220284
rect 307518 220084 307524 220148
rect 307588 220146 307594 220148
rect 316534 220146 316540 220148
rect 307588 220086 316540 220146
rect 307588 220084 307594 220086
rect 316534 220084 316540 220086
rect 316604 220084 316610 220148
rect 329230 220084 329236 220148
rect 329300 220146 329306 220148
rect 375966 220146 375972 220148
rect 329300 220086 375972 220146
rect 329300 220084 329306 220086
rect 375966 220084 375972 220086
rect 376036 220084 376042 220148
rect 324262 218996 324268 219060
rect 324332 219058 324338 219060
rect 336038 219058 336044 219060
rect 324332 218998 336044 219058
rect 324332 218996 324338 218998
rect 336038 218996 336044 218998
rect 336108 218996 336114 219060
rect 580758 218996 580764 219060
rect 580828 219058 580834 219060
rect 583520 219058 584960 219148
rect 580828 218998 584960 219058
rect 580828 218996 580834 218998
rect 326654 218860 326660 218924
rect 326724 218922 326730 218924
rect 358670 218922 358676 218924
rect 326724 218862 358676 218922
rect 326724 218860 326730 218862
rect 358670 218860 358676 218862
rect 358740 218860 358746 218924
rect 583520 218908 584960 218998
rect 319662 218724 319668 218788
rect 319732 218786 319738 218788
rect 353702 218786 353708 218788
rect 319732 218726 353708 218786
rect 319732 218724 319738 218726
rect 353702 218724 353708 218726
rect 353772 218724 353778 218788
rect 301998 218588 302004 218652
rect 302068 218650 302074 218652
rect 309910 218650 309916 218652
rect 302068 218590 309916 218650
rect 302068 218588 302074 218590
rect 309910 218588 309916 218590
rect 309980 218588 309986 218652
rect 311198 218588 311204 218652
rect 311268 218650 311274 218652
rect 327022 218650 327028 218652
rect 311268 218590 327028 218650
rect 311268 218588 311274 218590
rect 327022 218588 327028 218590
rect 327092 218588 327098 218652
rect 331070 218588 331076 218652
rect 331140 218650 331146 218652
rect 388478 218650 388484 218652
rect 331140 218590 388484 218650
rect 331140 218588 331146 218590
rect 388478 218588 388484 218590
rect 388548 218588 388554 218652
rect 318926 217500 318932 217564
rect 318996 217562 319002 217564
rect 351310 217562 351316 217564
rect 318996 217502 351316 217562
rect 318996 217500 319002 217502
rect 351310 217500 351316 217502
rect 351380 217500 351386 217564
rect 300526 217364 300532 217428
rect 300596 217426 300602 217428
rect 305126 217426 305132 217428
rect 300596 217366 305132 217426
rect 300596 217364 300602 217366
rect 305126 217364 305132 217366
rect 305196 217364 305202 217428
rect 319294 217364 319300 217428
rect 319364 217426 319370 217428
rect 352414 217426 352420 217428
rect 319364 217366 352420 217426
rect 319364 217364 319370 217366
rect 352414 217364 352420 217366
rect 352484 217364 352490 217428
rect 306782 217228 306788 217292
rect 306852 217290 306858 217292
rect 319478 217290 319484 217292
rect 306852 217230 319484 217290
rect 306852 217228 306858 217230
rect 319478 217228 319484 217230
rect 319548 217228 319554 217292
rect 329598 217228 329604 217292
rect 329668 217290 329674 217292
rect 378542 217290 378548 217292
rect 329668 217230 378548 217290
rect 329668 217228 329674 217230
rect 378542 217228 378548 217230
rect 378612 217228 378618 217292
rect 330702 217092 330708 217156
rect 330772 217154 330778 217156
rect 331990 217154 331996 217156
rect 330772 217094 331996 217154
rect 330772 217092 330778 217094
rect 331990 217092 331996 217094
rect 332060 217092 332066 217156
rect 325918 216684 325924 216748
rect 325988 216746 325994 216748
rect 329414 216746 329420 216748
rect 325988 216686 329420 216746
rect 325988 216684 325994 216686
rect 329414 216684 329420 216686
rect 329484 216684 329490 216748
rect 324446 216140 324452 216204
rect 324516 216202 324522 216204
rect 330518 216202 330524 216204
rect 324516 216142 330524 216202
rect 324516 216140 324522 216142
rect 330518 216140 330524 216142
rect 330588 216140 330594 216204
rect 332910 216140 332916 216204
rect 332980 216202 332986 216204
rect 338614 216202 338620 216204
rect 332980 216142 338620 216202
rect 332980 216140 332986 216142
rect 338614 216140 338620 216142
rect 338684 216140 338690 216204
rect 306414 216004 306420 216068
rect 306484 216066 306490 216068
rect 311014 216066 311020 216068
rect 306484 216006 311020 216066
rect 306484 216004 306490 216006
rect 311014 216004 311020 216006
rect 311084 216004 311090 216068
rect 314142 216004 314148 216068
rect 314212 216066 314218 216068
rect 324262 216066 324268 216068
rect 314212 216006 324268 216066
rect 314212 216004 314218 216006
rect 324262 216004 324268 216006
rect 324332 216004 324338 216068
rect 328310 216066 328316 216068
rect 325650 216006 328316 216066
rect 312670 215868 312676 215932
rect 312740 215930 312746 215932
rect 325650 215930 325710 216006
rect 328310 216004 328316 216006
rect 328380 216004 328386 216068
rect 328678 216004 328684 216068
rect 328748 216066 328754 216068
rect 360694 216066 360700 216068
rect 328748 216006 360700 216066
rect 328748 216004 328754 216006
rect 360694 216004 360700 216006
rect 360764 216004 360770 216068
rect 312740 215870 325710 215930
rect 312740 215868 312746 215870
rect 329966 215868 329972 215932
rect 330036 215930 330042 215932
rect 381118 215930 381124 215932
rect 330036 215870 381124 215930
rect 330036 215868 330042 215870
rect 381118 215868 381124 215870
rect 381188 215868 381194 215932
rect 327717 215794 327783 215797
rect 333094 215794 333100 215796
rect 327717 215792 333100 215794
rect 327717 215736 327722 215792
rect 327778 215736 333100 215792
rect 327717 215734 333100 215736
rect 327717 215731 327783 215734
rect 333094 215732 333100 215734
rect 333164 215732 333170 215796
rect 316350 215188 316356 215252
rect 316420 215250 316426 215252
rect 324998 215250 325004 215252
rect 316420 215190 325004 215250
rect 316420 215188 316426 215190
rect 324998 215188 325004 215190
rect 325068 215188 325074 215252
rect -960 214828 480 215068
rect 325182 214780 325188 214844
rect 325252 214842 325258 214844
rect 340086 214842 340092 214844
rect 325252 214782 340092 214842
rect 325252 214780 325258 214782
rect 340086 214780 340092 214782
rect 340156 214780 340162 214844
rect 332174 214644 332180 214708
rect 332244 214706 332250 214708
rect 356646 214706 356652 214708
rect 332244 214646 356652 214706
rect 332244 214644 332250 214646
rect 356646 214644 356652 214646
rect 356716 214644 356722 214708
rect 218973 214570 219039 214573
rect 281758 214570 281764 214572
rect 218973 214568 281764 214570
rect 218973 214512 218978 214568
rect 219034 214512 281764 214568
rect 218973 214510 281764 214512
rect 218973 214507 219039 214510
rect 281758 214508 281764 214510
rect 281828 214508 281834 214572
rect 312302 214508 312308 214572
rect 312372 214570 312378 214572
rect 330150 214570 330156 214572
rect 312372 214510 330156 214570
rect 312372 214508 312378 214510
rect 330150 214508 330156 214510
rect 330220 214508 330226 214572
rect 331806 214508 331812 214572
rect 331876 214570 331882 214572
rect 393630 214570 393636 214572
rect 331876 214510 393636 214570
rect 331876 214508 331882 214510
rect 393630 214508 393636 214510
rect 393700 214508 393706 214572
rect 302366 213964 302372 214028
rect 302436 214026 302442 214028
rect 310278 214026 310284 214028
rect 302436 213966 310284 214026
rect 302436 213964 302442 213966
rect 310278 213964 310284 213966
rect 310348 213964 310354 214028
rect 10174 213828 10180 213892
rect 10244 213890 10250 213892
rect 12382 213890 12388 213892
rect 10244 213830 12388 213890
rect 10244 213828 10250 213830
rect 12382 213828 12388 213830
rect 12452 213828 12458 213892
rect 1158 213148 1164 213212
rect 1228 213210 1234 213212
rect 11094 213210 11100 213212
rect 1228 213150 11100 213210
rect 1228 213148 1234 213150
rect 11094 213148 11100 213150
rect 11164 213148 11170 213212
rect 326470 213210 326476 213212
rect 322890 213150 326476 213210
rect 322890 213076 322950 213150
rect 326470 213148 326476 213150
rect 326540 213148 326546 213212
rect 311474 213012 311480 213076
rect 311544 213074 311550 213076
rect 312486 213074 312492 213076
rect 311544 213014 312492 213074
rect 311544 213012 311550 213014
rect 312486 213012 312492 213014
rect 312556 213012 312562 213076
rect 322882 213012 322888 213076
rect 322952 213012 322958 213076
rect 326194 213012 326200 213076
rect 326264 213074 326270 213076
rect 327574 213074 327580 213076
rect 326264 213014 327580 213074
rect 326264 213012 326270 213014
rect 327574 213012 327580 213014
rect 327644 213012 327650 213076
rect 328770 213012 328776 213076
rect 328840 213074 328846 213076
rect 334750 213074 334756 213076
rect 328840 213014 334756 213074
rect 328840 213012 328846 213014
rect 334750 213012 334756 213014
rect 334820 213012 334826 213076
rect 307753 212938 307819 212941
rect 327717 212940 327783 212941
rect 308530 212938 308536 212940
rect 307753 212936 308536 212938
rect 307753 212880 307758 212936
rect 307814 212880 308536 212936
rect 307753 212878 308536 212880
rect 307753 212875 307819 212878
rect 308530 212876 308536 212878
rect 308600 212876 308606 212940
rect 327666 212938 327672 212940
rect 327626 212878 327672 212938
rect 327736 212936 327783 212940
rect 327778 212880 327783 212936
rect 327666 212876 327672 212878
rect 327736 212876 327783 212880
rect 327717 212875 327783 212876
rect 583520 205580 584960 205820
rect -960 201922 480 202012
rect 2773 201922 2839 201925
rect -960 201920 2839 201922
rect -960 201864 2778 201920
rect 2834 201864 2839 201920
rect -960 201862 2839 201864
rect -960 201772 480 201862
rect 2773 201859 2839 201862
rect 281022 193156 281028 193220
rect 281092 193218 281098 193220
rect 284518 193218 284524 193220
rect 281092 193158 284524 193218
rect 281092 193156 281098 193158
rect 284518 193156 284524 193158
rect 284588 193156 284594 193220
rect 78438 192612 78444 192676
rect 78508 192674 78514 192676
rect 90030 192674 90036 192676
rect 78508 192614 90036 192674
rect 78508 192612 78514 192614
rect 90030 192612 90036 192614
rect 90100 192612 90106 192676
rect 89294 192476 89300 192540
rect 89364 192538 89370 192540
rect 110454 192538 110460 192540
rect 89364 192478 110460 192538
rect 89364 192476 89370 192478
rect 110454 192476 110460 192478
rect 110524 192476 110530 192540
rect 283833 192538 283899 192541
rect 290457 192538 290523 192541
rect 283833 192536 290523 192538
rect 283833 192480 283838 192536
rect 283894 192480 290462 192536
rect 290518 192480 290523 192536
rect 283833 192478 290523 192480
rect 283833 192475 283899 192478
rect 290457 192475 290523 192478
rect 580901 192538 580967 192541
rect 583520 192538 584960 192628
rect 580901 192536 584960 192538
rect 580901 192480 580906 192536
rect 580962 192480 584960 192536
rect 580901 192478 584960 192480
rect 580901 192475 580967 192478
rect 583520 192388 584960 192478
rect 287053 191994 287119 191997
rect 298093 191994 298159 191997
rect 287053 191992 298159 191994
rect 287053 191936 287058 191992
rect 287114 191936 298098 191992
rect 298154 191936 298159 191992
rect 287053 191934 298159 191936
rect 287053 191931 287119 191934
rect 298093 191931 298159 191934
rect 281809 191858 281875 191861
rect 301078 191858 301084 191860
rect 281809 191856 301084 191858
rect 281809 191800 281814 191856
rect 281870 191800 301084 191856
rect 281809 191798 301084 191800
rect 281809 191795 281875 191798
rect 301078 191796 301084 191798
rect 301148 191796 301154 191860
rect 335118 191796 335124 191860
rect 335188 191858 335194 191860
rect 337326 191858 337332 191860
rect 335188 191798 337332 191858
rect 335188 191796 335194 191798
rect 337326 191796 337332 191798
rect 337396 191796 337402 191860
rect 2630 190980 2636 191044
rect 2700 191042 2706 191044
rect 10174 191042 10180 191044
rect 2700 190982 10180 191042
rect 2700 190980 2706 190982
rect 10174 190980 10180 190982
rect 10244 190980 10250 191044
rect 281901 190770 281967 190773
rect 298686 190770 298692 190772
rect 281901 190768 298692 190770
rect 281901 190712 281906 190768
rect 281962 190712 298692 190768
rect 281901 190710 298692 190712
rect 281901 190707 281967 190710
rect 298686 190708 298692 190710
rect 298756 190708 298762 190772
rect 281390 190572 281396 190636
rect 281460 190634 281466 190636
rect 300485 190634 300551 190637
rect 281460 190632 300551 190634
rect 281460 190576 300490 190632
rect 300546 190576 300551 190632
rect 281460 190574 300551 190576
rect 281460 190572 281466 190574
rect 300485 190571 300551 190574
rect 282862 190436 282868 190500
rect 282932 190498 282938 190500
rect 291694 190498 291700 190500
rect 282932 190438 291700 190498
rect 282932 190436 282938 190438
rect 291694 190436 291700 190438
rect 291764 190436 291770 190500
rect 298686 190436 298692 190500
rect 298756 190498 298762 190500
rect 302325 190498 302391 190501
rect 298756 190496 302391 190498
rect 298756 190440 302330 190496
rect 302386 190440 302391 190496
rect 298756 190438 302391 190440
rect 298756 190436 298762 190438
rect 302325 190435 302391 190438
rect 9622 190300 9628 190364
rect 9692 190362 9698 190364
rect 9857 190362 9923 190365
rect 9692 190360 9923 190362
rect 9692 190304 9862 190360
rect 9918 190304 9923 190360
rect 9692 190302 9923 190304
rect 9692 190300 9698 190302
rect 9857 190299 9923 190302
rect 283782 189620 283788 189684
rect 283852 189682 283858 189684
rect 299790 189682 299796 189684
rect 283852 189622 299796 189682
rect 283852 189620 283858 189622
rect 299790 189620 299796 189622
rect 299860 189620 299866 189684
rect 283046 189484 283052 189548
rect 283116 189546 283122 189548
rect 300945 189546 301011 189549
rect 283116 189544 301011 189546
rect 283116 189488 300950 189544
rect 301006 189488 301011 189544
rect 283116 189486 301011 189488
rect 283116 189484 283122 189486
rect 300945 189483 301011 189486
rect 284293 189410 284359 189413
rect 299974 189410 299980 189412
rect 284293 189408 299980 189410
rect 284293 189352 284298 189408
rect 284354 189352 299980 189408
rect 284293 189350 299980 189352
rect 284293 189347 284359 189350
rect 299974 189348 299980 189350
rect 300044 189348 300050 189412
rect 282494 189212 282500 189276
rect 282564 189274 282570 189276
rect 292798 189274 292804 189276
rect 282564 189214 292804 189274
rect 282564 189212 282570 189214
rect 292798 189212 292804 189214
rect 292868 189212 292874 189276
rect 300485 189274 300551 189277
rect 302233 189274 302299 189277
rect 300485 189272 302299 189274
rect 300485 189216 300490 189272
rect 300546 189216 302238 189272
rect 302294 189216 302299 189272
rect 300485 189214 302299 189216
rect 300485 189211 300551 189214
rect 302233 189211 302299 189214
rect 281612 189078 281826 189138
rect 281766 189002 281826 189078
rect 283966 189076 283972 189140
rect 284036 189138 284042 189140
rect 297541 189138 297607 189141
rect 284036 189136 297607 189138
rect 284036 189080 297546 189136
rect 297602 189080 297607 189136
rect 284036 189078 297607 189080
rect 284036 189076 284042 189078
rect 297541 189075 297607 189078
rect 302374 189078 302588 189138
rect -960 188866 480 188956
rect 281704 188942 281826 189002
rect 2773 188866 2839 188869
rect 281766 188866 281826 188942
rect -960 188864 2839 188866
rect -960 188808 2778 188864
rect 2834 188808 2839 188864
rect -960 188806 2839 188808
rect 281612 188806 281826 188866
rect -960 188716 480 188806
rect 2773 188803 2839 188806
rect 281674 188730 281734 188806
rect 281612 188670 281734 188730
rect 281674 188594 281734 188670
rect 285806 188668 285812 188732
rect 285876 188730 285882 188732
rect 301262 188730 301268 188732
rect 285876 188670 301268 188730
rect 285876 188668 285882 188670
rect 301262 188668 301268 188670
rect 301332 188668 301338 188732
rect 281612 188534 281826 188594
rect 281766 188322 281826 188534
rect 284150 188532 284156 188596
rect 284220 188594 284226 188596
rect 296846 188594 296852 188596
rect 284220 188534 296852 188594
rect 284220 188532 284226 188534
rect 296846 188532 296852 188534
rect 296916 188532 296922 188596
rect 302374 188458 302434 189078
rect 302740 189004 302804 189010
rect 302740 188934 302804 188940
rect 302734 188804 302740 188868
rect 302804 188866 302810 188868
rect 302804 188806 303630 188866
rect 302804 188804 302810 188806
rect 303570 188730 303630 188806
rect 303508 188670 303630 188730
rect 303570 188594 303630 188670
rect 303508 188534 303630 188594
rect 302374 188398 302588 188458
rect 281612 188262 281826 188322
rect 292982 188260 292988 188324
rect 293052 188322 293058 188324
rect 300894 188322 300900 188324
rect 293052 188262 300900 188322
rect 293052 188260 293058 188262
rect 300894 188260 300900 188262
rect 300964 188260 300970 188324
rect 302734 188260 302740 188324
rect 302804 188260 302810 188324
rect 302464 188188 302528 188194
rect 281704 188126 302464 188186
rect 302464 188118 302528 188124
rect 291142 188050 291148 188052
rect 281612 187990 291148 188050
rect 291142 187988 291148 187990
rect 291212 188050 291218 188052
rect 291212 187990 302588 188050
rect 291212 187988 291218 187990
rect 281809 187914 281875 187917
rect 281612 187912 281875 187914
rect 281612 187856 281814 187912
rect 281870 187856 281875 187912
rect 281612 187854 281875 187856
rect 281809 187851 281875 187854
rect 283414 187852 283420 187916
rect 283484 187914 283490 187916
rect 292614 187914 292620 187916
rect 283484 187854 292620 187914
rect 283484 187852 283490 187854
rect 292614 187852 292620 187854
rect 292684 187852 292690 187916
rect 301078 187852 301084 187916
rect 301148 187914 301154 187916
rect 301446 187914 301452 187916
rect 301148 187854 301452 187914
rect 301148 187852 301154 187854
rect 301446 187852 301452 187854
rect 301516 187914 301522 187916
rect 301516 187854 302588 187914
rect 301516 187852 301522 187854
rect 295977 187778 296043 187781
rect 281612 187776 302588 187778
rect 281612 187720 295982 187776
rect 296038 187720 302588 187776
rect 281612 187718 302588 187720
rect 295977 187715 296043 187718
rect 299238 187642 299244 187644
rect 281704 187582 299244 187642
rect 299238 187580 299244 187582
rect 299308 187642 299314 187644
rect 299308 187582 302496 187642
rect 299308 187580 299314 187582
rect 284293 187506 284359 187509
rect 281704 187504 284359 187506
rect 281704 187448 284298 187504
rect 284354 187448 284359 187504
rect 281704 187446 284359 187448
rect 284293 187443 284359 187446
rect 299974 187444 299980 187508
rect 300044 187506 300050 187508
rect 300044 187446 302496 187506
rect 300044 187444 300050 187446
rect 281390 187308 281396 187372
rect 281460 187308 281466 187372
rect 302233 187370 302299 187373
rect 302233 187368 302588 187370
rect 302233 187312 302238 187368
rect 302294 187312 302588 187368
rect 302233 187310 302588 187312
rect 302233 187307 302299 187310
rect 283782 187234 283788 187236
rect 281612 187174 283788 187234
rect 283782 187172 283788 187174
rect 283852 187172 283858 187236
rect 299790 187172 299796 187236
rect 299860 187234 299866 187236
rect 300158 187234 300164 187236
rect 299860 187174 300164 187234
rect 299860 187172 299866 187174
rect 300158 187172 300164 187174
rect 300228 187234 300234 187236
rect 300228 187174 302588 187234
rect 300228 187172 300234 187174
rect 300710 187098 300716 187100
rect 281612 187038 300716 187098
rect 300710 187036 300716 187038
rect 300780 187098 300786 187100
rect 300780 187038 302588 187098
rect 300780 187036 300786 187038
rect 298185 186962 298251 186965
rect 281612 186960 302588 186962
rect 281612 186904 298190 186960
rect 298246 186904 302588 186960
rect 281612 186902 302588 186904
rect 298185 186899 298251 186902
rect 281809 186826 281875 186829
rect 281612 186824 281875 186826
rect 281612 186768 281814 186824
rect 281870 186768 281875 186824
rect 281612 186766 281875 186768
rect 281809 186763 281875 186766
rect 284334 186764 284340 186828
rect 284404 186826 284410 186828
rect 285581 186826 285647 186829
rect 284404 186824 285647 186826
rect 284404 186768 285586 186824
rect 285642 186768 285647 186824
rect 284404 186766 285647 186768
rect 284404 186764 284410 186766
rect 285581 186763 285647 186766
rect 291837 186826 291903 186829
rect 297950 186826 297956 186828
rect 291837 186824 297956 186826
rect 291837 186768 291842 186824
rect 291898 186768 297956 186824
rect 291837 186766 297956 186768
rect 291837 186763 291903 186766
rect 297950 186764 297956 186766
rect 298020 186764 298026 186828
rect 298093 186826 298159 186829
rect 298093 186824 302588 186826
rect 298093 186768 298098 186824
rect 298154 186768 302588 186824
rect 298093 186766 302588 186768
rect 298093 186763 298159 186766
rect 281901 186690 281967 186693
rect 281612 186688 281967 186690
rect 281612 186632 281906 186688
rect 281962 186632 281967 186688
rect 281612 186630 281967 186632
rect 281901 186627 281967 186630
rect 283598 186628 283604 186692
rect 283668 186690 283674 186692
rect 297398 186690 297404 186692
rect 283668 186630 297404 186690
rect 283668 186628 283674 186630
rect 297398 186628 297404 186630
rect 297468 186690 297474 186692
rect 299422 186690 299428 186692
rect 297468 186630 299428 186690
rect 297468 186628 297474 186630
rect 299422 186628 299428 186630
rect 299492 186628 299498 186692
rect 302325 186690 302391 186693
rect 302325 186688 302588 186690
rect 302325 186632 302330 186688
rect 302386 186632 302588 186688
rect 302325 186630 302588 186632
rect 302325 186627 302391 186630
rect 298134 186554 298140 186556
rect 281612 186494 298140 186554
rect 298134 186492 298140 186494
rect 298204 186554 298210 186556
rect 298204 186494 302588 186554
rect 298204 186492 298210 186494
rect 291837 186418 291903 186421
rect 281612 186416 291903 186418
rect 281612 186360 291842 186416
rect 291898 186360 291903 186416
rect 281612 186358 291903 186360
rect 291837 186355 291903 186358
rect 297950 186356 297956 186420
rect 298020 186418 298026 186420
rect 298020 186358 302588 186418
rect 298020 186356 298026 186358
rect 283598 186282 283604 186284
rect 281612 186222 283604 186282
rect 283598 186220 283604 186222
rect 283668 186220 283674 186284
rect 299422 186220 299428 186284
rect 299492 186282 299498 186284
rect 299492 186222 302588 186282
rect 299492 186220 299498 186222
rect 283966 186146 283972 186148
rect 281704 186086 283972 186146
rect 283966 186084 283972 186086
rect 284036 186084 284042 186148
rect 297541 186146 297607 186149
rect 297541 186144 302496 186146
rect 297541 186088 297546 186144
rect 297602 186088 302496 186144
rect 297541 186086 302496 186088
rect 297541 186083 297607 186086
rect 284150 186010 284156 186012
rect 281612 185950 284156 186010
rect 284150 185948 284156 185950
rect 284220 185948 284226 186012
rect 296846 185948 296852 186012
rect 296916 186010 296922 186012
rect 296916 185950 302588 186010
rect 296916 185948 296922 185950
rect 296294 185874 296300 185876
rect 281612 185814 296300 185874
rect 296294 185812 296300 185814
rect 296364 185812 296370 185876
rect 299790 185812 299796 185876
rect 299860 185874 299866 185876
rect 299860 185814 302588 185874
rect 299860 185812 299866 185814
rect 295926 185738 295932 185740
rect 281612 185678 295932 185738
rect 295926 185676 295932 185678
rect 295996 185738 296002 185740
rect 295996 185678 302588 185738
rect 295996 185676 296002 185678
rect 295558 185602 295564 185604
rect 281612 185542 295564 185602
rect 295558 185540 295564 185542
rect 295628 185602 295634 185604
rect 295628 185542 302588 185602
rect 295628 185540 295634 185542
rect 295190 185466 295196 185468
rect 281612 185406 295196 185466
rect 295190 185404 295196 185406
rect 295260 185466 295266 185468
rect 295260 185406 302588 185466
rect 295260 185404 295266 185406
rect 294822 185330 294828 185332
rect 281612 185270 294828 185330
rect 294822 185268 294828 185270
rect 294892 185330 294898 185332
rect 294892 185270 302588 185330
rect 294892 185268 294898 185270
rect 294454 185194 294460 185196
rect 281612 185134 294460 185194
rect 294454 185132 294460 185134
rect 294524 185194 294530 185196
rect 294524 185134 302588 185194
rect 294524 185132 294530 185134
rect 294086 185058 294092 185060
rect 281612 184998 294092 185058
rect 294086 184996 294092 184998
rect 294156 185058 294162 185060
rect 294156 184998 302588 185058
rect 294156 184996 294162 184998
rect 283414 184922 283420 184924
rect 281612 184862 283420 184922
rect 283414 184860 283420 184862
rect 283484 184860 283490 184924
rect 287094 184860 287100 184924
rect 287164 184922 287170 184924
rect 288341 184922 288407 184925
rect 287164 184920 288407 184922
rect 287164 184864 288346 184920
rect 288402 184864 288407 184920
rect 287164 184862 288407 184864
rect 287164 184860 287170 184862
rect 288341 184859 288407 184862
rect 292614 184860 292620 184924
rect 292684 184922 292690 184924
rect 293718 184922 293724 184924
rect 292684 184862 293724 184922
rect 292684 184860 292690 184862
rect 293718 184860 293724 184862
rect 293788 184922 293794 184924
rect 293788 184862 302588 184922
rect 293788 184860 293794 184862
rect 282494 184786 282500 184788
rect 281612 184726 282500 184786
rect 282494 184724 282500 184726
rect 282564 184724 282570 184788
rect 282913 184786 282979 184789
rect 284201 184786 284267 184789
rect 287053 184786 287119 184789
rect 282913 184784 287119 184786
rect 282913 184728 282918 184784
rect 282974 184728 284206 184784
rect 284262 184728 287058 184784
rect 287114 184728 287119 184784
rect 282913 184726 287119 184728
rect 282913 184723 282979 184726
rect 284201 184723 284267 184726
rect 287053 184723 287119 184726
rect 292798 184724 292804 184788
rect 292868 184786 292874 184788
rect 293350 184786 293356 184788
rect 292868 184726 293356 184786
rect 292868 184724 292874 184726
rect 293350 184724 293356 184726
rect 293420 184786 293426 184788
rect 293420 184726 302588 184786
rect 293420 184724 293426 184726
rect 282126 184650 282132 184652
rect 281612 184590 282132 184650
rect 282126 184588 282132 184590
rect 282196 184588 282202 184652
rect 299974 184588 299980 184652
rect 300044 184650 300050 184652
rect 300761 184650 300827 184653
rect 300044 184648 300827 184650
rect 300044 184592 300766 184648
rect 300822 184592 300827 184648
rect 300044 184590 300827 184592
rect 300044 184588 300050 184590
rect 300761 184587 300827 184590
rect 300894 184588 300900 184652
rect 300964 184650 300970 184652
rect 300964 184590 302588 184650
rect 300964 184588 300970 184590
rect 292614 184514 292620 184516
rect 281612 184454 292620 184514
rect 292614 184452 292620 184454
rect 292684 184514 292690 184516
rect 292684 184454 302588 184514
rect 292684 184452 292690 184454
rect 282678 184378 282684 184380
rect 281612 184318 282684 184378
rect 282678 184316 282684 184318
rect 282748 184316 282754 184380
rect 301630 184316 301636 184380
rect 301700 184378 301706 184380
rect 301700 184318 302588 184378
rect 301700 184316 301706 184318
rect 281809 184242 281875 184245
rect 281612 184240 281875 184242
rect 281612 184184 281814 184240
rect 281870 184184 281875 184240
rect 281612 184182 281875 184184
rect 281809 184179 281875 184182
rect 299565 184242 299631 184245
rect 299565 184240 302588 184242
rect 299565 184184 299570 184240
rect 299626 184184 302588 184240
rect 299565 184182 302588 184184
rect 299565 184179 299631 184182
rect 291510 184106 291516 184108
rect 281704 184046 291516 184106
rect 291510 184044 291516 184046
rect 291580 184106 291586 184108
rect 291580 184046 302496 184106
rect 291580 184044 291586 184046
rect 290222 183970 290228 183972
rect 281612 183910 290228 183970
rect 290222 183908 290228 183910
rect 290292 183970 290298 183972
rect 290292 183910 302588 183970
rect 290292 183908 290298 183910
rect 291837 183836 291903 183837
rect 290590 183834 290596 183836
rect 281612 183774 290596 183834
rect 290590 183772 290596 183774
rect 290660 183772 290666 183836
rect 291837 183832 291884 183836
rect 291948 183834 291954 183836
rect 299565 183834 299631 183837
rect 291948 183832 299631 183834
rect 291837 183776 291842 183832
rect 291948 183776 299570 183832
rect 299626 183776 299631 183832
rect 291837 183772 291884 183776
rect 291948 183774 299631 183776
rect 291948 183772 291954 183774
rect 291837 183771 291903 183772
rect 299565 183771 299631 183774
rect 300526 183772 300532 183836
rect 300596 183834 300602 183836
rect 300596 183774 302588 183834
rect 300596 183772 300602 183774
rect 289486 183698 289492 183700
rect 281612 183638 289492 183698
rect 289486 183636 289492 183638
rect 289556 183698 289562 183700
rect 289556 183638 302588 183698
rect 289556 183636 289562 183638
rect 284109 183562 284175 183565
rect 281612 183560 284175 183562
rect 281612 183504 284114 183560
rect 284170 183504 284175 183560
rect 281612 183502 284175 183504
rect 284109 183499 284175 183502
rect 289670 183500 289676 183564
rect 289740 183562 289746 183564
rect 289740 183502 302588 183562
rect 289740 183500 289746 183502
rect 288934 183426 288940 183428
rect 281704 183366 288940 183426
rect 288934 183364 288940 183366
rect 289004 183426 289010 183428
rect 289004 183366 302496 183426
rect 289004 183364 289010 183366
rect 282821 183290 282887 183293
rect 281612 183288 282887 183290
rect 281612 183232 282826 183288
rect 282882 183232 282887 183288
rect 281612 183230 282887 183232
rect 282821 183227 282887 183230
rect 284109 183290 284175 183293
rect 289302 183290 289308 183292
rect 284109 183288 289308 183290
rect 284109 183232 284114 183288
rect 284170 183232 289308 183288
rect 284109 183230 289308 183232
rect 284109 183227 284175 183230
rect 289302 183228 289308 183230
rect 289372 183290 289378 183292
rect 289670 183290 289676 183292
rect 289372 183230 289676 183290
rect 289372 183228 289378 183230
rect 289670 183228 289676 183230
rect 289740 183228 289746 183292
rect 300853 183290 300919 183293
rect 300853 183288 302588 183290
rect 300853 183232 300858 183288
rect 300914 183232 302588 183288
rect 300853 183230 302588 183232
rect 300853 183227 300919 183230
rect 288198 183154 288204 183156
rect 281704 183094 288204 183154
rect 288198 183092 288204 183094
rect 288268 183154 288274 183156
rect 288268 183094 302496 183154
rect 288268 183092 288274 183094
rect 287830 183018 287836 183020
rect 281612 182958 287836 183018
rect 287830 182956 287836 182958
rect 287900 183018 287906 183020
rect 287900 182958 302588 183018
rect 287900 182956 287906 182958
rect 287462 182882 287468 182884
rect 281612 182822 287468 182882
rect 287462 182820 287468 182822
rect 287532 182882 287538 182884
rect 287532 182822 302588 182882
rect 287532 182820 287538 182822
rect 287094 182746 287100 182748
rect 281612 182686 287100 182746
rect 287094 182684 287100 182686
rect 287164 182746 287170 182748
rect 287164 182686 302588 182746
rect 287164 182684 287170 182686
rect 281809 182610 281875 182613
rect 281612 182608 281875 182610
rect 281612 182552 281814 182608
rect 281870 182552 281875 182608
rect 281612 182550 281875 182552
rect 281809 182547 281875 182550
rect 301078 182548 301084 182612
rect 301148 182610 301154 182612
rect 301148 182550 302588 182610
rect 301148 182548 301154 182550
rect 281022 182412 281028 182476
rect 281092 182412 281098 182476
rect 300894 182412 300900 182476
rect 300964 182474 300970 182476
rect 300964 182414 302588 182474
rect 300964 182412 300970 182414
rect 285990 182338 285996 182340
rect 281612 182278 285996 182338
rect 285990 182276 285996 182278
rect 286060 182338 286066 182340
rect 286060 182278 302588 182338
rect 286060 182276 286066 182278
rect 288617 182204 288683 182205
rect 285806 182202 285812 182204
rect 281612 182142 285812 182202
rect 285806 182140 285812 182142
rect 285876 182140 285882 182204
rect 288566 182202 288572 182204
rect 288526 182142 288572 182202
rect 288636 182200 288683 182204
rect 288678 182144 288683 182200
rect 288566 182140 288572 182142
rect 288636 182140 288683 182144
rect 301262 182140 301268 182204
rect 301332 182202 301338 182204
rect 301332 182142 302588 182202
rect 301332 182140 301338 182142
rect 288617 182139 288683 182140
rect 285254 182066 285260 182068
rect 281612 182006 285260 182066
rect 285254 182004 285260 182006
rect 285324 182066 285330 182068
rect 285324 182006 302588 182066
rect 285324 182004 285330 182006
rect 281901 181930 281967 181933
rect 281612 181928 281967 181930
rect 281612 181872 281906 181928
rect 281962 181872 281967 181928
rect 281612 181870 281967 181872
rect 281901 181867 281967 181870
rect 302233 181930 302299 181933
rect 302233 181928 302588 181930
rect 302233 181872 302238 181928
rect 302294 181872 302588 181928
rect 302233 181870 302588 181872
rect 302233 181867 302299 181870
rect 285438 181794 285444 181796
rect 281612 181734 285444 181794
rect 285438 181732 285444 181734
rect 285508 181794 285514 181796
rect 285508 181734 302588 181794
rect 285508 181732 285514 181734
rect 281574 181596 281580 181660
rect 281644 181658 281650 181660
rect 281644 181598 302588 181658
rect 281644 181596 281650 181598
rect 284150 181522 284156 181524
rect 281704 181462 284156 181522
rect 284150 181460 284156 181462
rect 284220 181522 284226 181524
rect 284220 181462 302496 181522
rect 284220 181460 284226 181462
rect 281809 181386 281875 181389
rect 283046 181386 283052 181388
rect 281612 181384 283052 181386
rect 281612 181328 281814 181384
rect 281870 181328 283052 181384
rect 281612 181326 283052 181328
rect 281809 181323 281875 181326
rect 283046 181324 283052 181326
rect 283116 181324 283122 181388
rect 300945 181386 301011 181389
rect 300945 181384 302588 181386
rect 300945 181328 300950 181384
rect 301006 181328 302588 181384
rect 300945 181326 302588 181328
rect 300945 181323 301011 181326
rect 283046 181250 283052 181252
rect 281612 181190 283052 181250
rect 283046 181188 283052 181190
rect 283116 181250 283122 181252
rect 283116 181190 302588 181250
rect 283116 181188 283122 181190
rect 284702 181114 284708 181116
rect 281704 181054 284708 181114
rect 284702 181052 284708 181054
rect 284772 181114 284778 181116
rect 284772 181054 302496 181114
rect 284772 181052 284778 181054
rect 281390 180916 281396 180980
rect 281460 180916 281466 180980
rect 302182 180916 302188 180980
rect 302252 180978 302258 180980
rect 302252 180918 302588 180978
rect 302252 180916 302258 180918
rect 282678 180842 282684 180844
rect 281612 180782 282684 180842
rect 282678 180780 282684 180782
rect 282748 180842 282754 180844
rect 282748 180782 302588 180842
rect 282748 180780 282754 180782
rect 281574 180644 281580 180708
rect 281644 180706 281650 180708
rect 281644 180646 302588 180706
rect 281644 180644 281650 180646
rect 281582 180434 281642 180540
rect 281950 180510 302496 180570
rect 281950 180434 282010 180510
rect 281582 180374 282010 180434
rect 281582 180029 281642 180374
rect 282126 180372 282132 180436
rect 282196 180434 282202 180436
rect 292982 180434 292988 180436
rect 282196 180374 292988 180434
rect 282196 180372 282202 180374
rect 292982 180372 292988 180374
rect 293052 180372 293058 180436
rect 296621 180434 296687 180437
rect 296846 180434 296852 180436
rect 296576 180432 296852 180434
rect 296576 180376 296626 180432
rect 296682 180376 296852 180432
rect 296576 180374 296852 180376
rect 296621 180371 296687 180374
rect 296846 180372 296852 180374
rect 296916 180372 296922 180436
rect 290590 180236 290596 180300
rect 290660 180298 290666 180300
rect 300526 180298 300532 180300
rect 290660 180238 300532 180298
rect 290660 180236 290666 180238
rect 300526 180236 300532 180238
rect 300596 180236 300602 180300
rect 288341 180162 288407 180165
rect 300158 180162 300164 180164
rect 288341 180160 300164 180162
rect 288341 180104 288346 180160
rect 288402 180104 300164 180160
rect 288341 180102 300164 180104
rect 288341 180099 288407 180102
rect 300158 180100 300164 180102
rect 300228 180100 300234 180164
rect 281582 180024 281691 180029
rect 281582 179968 281630 180024
rect 281686 179968 281691 180024
rect 281582 179966 281691 179968
rect 281625 179963 281691 179966
rect 285581 180026 285647 180029
rect 285581 180024 296730 180026
rect 285581 179968 285586 180024
rect 285642 179968 296730 180024
rect 285581 179966 296730 179968
rect 285581 179963 285647 179966
rect 296670 179890 296730 179966
rect 302550 179890 302556 179892
rect 296670 179830 302556 179890
rect 302550 179828 302556 179830
rect 302620 179828 302626 179892
rect 298870 179692 298876 179756
rect 298940 179754 298946 179756
rect 300894 179754 300900 179756
rect 298940 179694 300900 179754
rect 298940 179692 298946 179694
rect 300894 179692 300900 179694
rect 300964 179692 300970 179756
rect 299238 179556 299244 179620
rect 299308 179618 299314 179620
rect 302233 179618 302299 179621
rect 299308 179616 302299 179618
rect 299308 179560 302238 179616
rect 302294 179560 302299 179616
rect 299308 179558 302299 179560
rect 299308 179556 299314 179558
rect 302233 179555 302299 179558
rect 290038 179420 290044 179484
rect 290108 179482 290114 179484
rect 290590 179482 290596 179484
rect 290108 179422 290596 179482
rect 290108 179420 290114 179422
rect 290590 179420 290596 179422
rect 290660 179420 290666 179484
rect 300761 179482 300827 179485
rect 301497 179482 301563 179485
rect 300761 179480 301563 179482
rect 300761 179424 300766 179480
rect 300822 179424 301502 179480
rect 301558 179424 301563 179480
rect 300761 179422 301563 179424
rect 300761 179419 300827 179422
rect 301497 179419 301563 179422
rect 182122 179284 182128 179348
rect 182192 179346 182198 179348
rect 182858 179346 182864 179348
rect 182192 179286 182864 179346
rect 182192 179284 182198 179286
rect 182858 179284 182864 179286
rect 182928 179346 182934 179348
rect 183594 179346 183600 179348
rect 182928 179286 183600 179346
rect 182928 179284 182934 179286
rect 183594 179284 183600 179286
rect 183664 179346 183670 179348
rect 184330 179346 184336 179348
rect 183664 179286 184336 179346
rect 183664 179284 183670 179286
rect 184330 179284 184336 179286
rect 184400 179346 184406 179348
rect 185066 179346 185072 179348
rect 184400 179286 185072 179346
rect 184400 179284 184406 179286
rect 185066 179284 185072 179286
rect 185136 179346 185142 179348
rect 186538 179346 186544 179348
rect 185136 179286 186544 179346
rect 185136 179284 185142 179286
rect 185810 179212 185870 179286
rect 186538 179284 186544 179286
rect 186608 179346 186614 179348
rect 187274 179346 187280 179348
rect 186608 179286 187280 179346
rect 186608 179284 186614 179286
rect 187274 179284 187280 179286
rect 187344 179346 187350 179348
rect 188010 179346 188016 179348
rect 187344 179286 188016 179346
rect 187344 179284 187350 179286
rect 188010 179284 188016 179286
rect 188080 179346 188086 179348
rect 188746 179346 188752 179348
rect 188080 179286 188752 179346
rect 188080 179284 188086 179286
rect 188746 179284 188752 179286
rect 188816 179346 188822 179348
rect 189482 179346 189488 179348
rect 188816 179286 189488 179346
rect 188816 179284 188822 179286
rect 189482 179284 189488 179286
rect 189552 179346 189558 179348
rect 190218 179346 190224 179348
rect 189552 179286 190224 179346
rect 189552 179284 189558 179286
rect 190218 179284 190224 179286
rect 190288 179346 190294 179348
rect 191690 179346 191696 179348
rect 190288 179286 191696 179346
rect 190288 179284 190294 179286
rect 190962 179212 191022 179286
rect 191690 179284 191696 179286
rect 191760 179346 191766 179348
rect 192426 179346 192432 179348
rect 191760 179286 192432 179346
rect 191760 179284 191766 179286
rect 192426 179284 192432 179286
rect 192496 179346 192502 179348
rect 193162 179346 193168 179348
rect 192496 179286 193168 179346
rect 192496 179284 192502 179286
rect 193162 179284 193168 179286
rect 193232 179346 193238 179348
rect 193898 179346 193904 179348
rect 193232 179286 193904 179346
rect 193232 179284 193238 179286
rect 193898 179284 193904 179286
rect 193968 179346 193974 179348
rect 194634 179346 194640 179348
rect 193968 179286 194640 179346
rect 193968 179284 193974 179286
rect 194634 179284 194640 179286
rect 194704 179346 194710 179348
rect 195370 179346 195376 179348
rect 194704 179286 195376 179346
rect 194704 179284 194710 179286
rect 195370 179284 195376 179286
rect 195440 179346 195446 179348
rect 196106 179346 196112 179348
rect 195440 179286 196112 179346
rect 195440 179284 195446 179286
rect 196106 179284 196112 179286
rect 196176 179346 196182 179348
rect 196842 179346 196848 179348
rect 196176 179286 196848 179346
rect 196176 179284 196182 179286
rect 196842 179284 196848 179286
rect 196912 179346 196918 179348
rect 197578 179346 197584 179348
rect 196912 179286 197584 179346
rect 196912 179284 196918 179286
rect 197578 179284 197584 179286
rect 197648 179346 197654 179348
rect 198314 179346 198320 179348
rect 197648 179286 198320 179346
rect 197648 179284 197654 179286
rect 198314 179284 198320 179286
rect 198384 179284 198390 179348
rect 214782 179284 214788 179348
rect 214852 179346 214858 179348
rect 215518 179346 215524 179348
rect 214852 179286 215524 179346
rect 214852 179284 214858 179286
rect 215518 179284 215524 179286
rect 215588 179346 215594 179348
rect 216254 179346 216260 179348
rect 215588 179286 216260 179346
rect 215588 179284 215594 179286
rect 216254 179284 216260 179286
rect 216324 179346 216330 179348
rect 216990 179346 216996 179348
rect 216324 179286 216996 179346
rect 216324 179284 216330 179286
rect 216990 179284 216996 179286
rect 217060 179346 217066 179348
rect 217726 179346 217732 179348
rect 217060 179286 217732 179346
rect 217060 179284 217066 179286
rect 217726 179284 217732 179286
rect 217796 179346 217802 179348
rect 218462 179346 218468 179348
rect 217796 179286 218468 179346
rect 217796 179284 217802 179286
rect 218462 179284 218468 179286
rect 218532 179346 218538 179348
rect 219198 179346 219204 179348
rect 218532 179286 219204 179346
rect 218532 179284 218538 179286
rect 219198 179284 219204 179286
rect 219268 179346 219274 179348
rect 219934 179346 219940 179348
rect 219268 179286 219940 179346
rect 219268 179284 219274 179286
rect 219934 179284 219940 179286
rect 220004 179346 220010 179348
rect 220854 179346 220860 179348
rect 220004 179286 220860 179346
rect 220004 179284 220010 179286
rect 220854 179284 220860 179286
rect 220924 179346 220930 179348
rect 221406 179346 221412 179348
rect 220924 179286 221412 179346
rect 220924 179284 220930 179286
rect 221406 179284 221412 179286
rect 221476 179346 221482 179348
rect 222142 179346 222148 179348
rect 221476 179286 222148 179346
rect 221476 179284 221482 179286
rect 222142 179284 222148 179286
rect 222212 179346 222218 179348
rect 222878 179346 222884 179348
rect 222212 179286 222884 179346
rect 222212 179284 222218 179286
rect 222878 179284 222884 179286
rect 222948 179346 222954 179348
rect 223614 179346 223620 179348
rect 222948 179286 223620 179346
rect 222948 179284 222954 179286
rect 223614 179284 223620 179286
rect 223684 179284 223690 179348
rect 248914 179284 248920 179348
rect 248984 179346 248990 179348
rect 249650 179346 249656 179348
rect 248984 179286 249656 179346
rect 248984 179284 248990 179286
rect 249650 179284 249656 179286
rect 249720 179346 249726 179348
rect 250386 179346 250392 179348
rect 249720 179286 250392 179346
rect 249720 179284 249726 179286
rect 250386 179284 250392 179286
rect 250456 179346 250462 179348
rect 251122 179346 251128 179348
rect 250456 179286 251128 179346
rect 250456 179284 250462 179286
rect 251122 179284 251128 179286
rect 251192 179346 251198 179348
rect 251858 179346 251864 179348
rect 251192 179286 251864 179346
rect 251192 179284 251198 179286
rect 251858 179284 251864 179286
rect 251928 179346 251934 179348
rect 252594 179346 252600 179348
rect 251928 179286 252600 179346
rect 251928 179284 251934 179286
rect 252594 179284 252600 179286
rect 252664 179346 252670 179348
rect 253330 179346 253336 179348
rect 252664 179286 253336 179346
rect 252664 179284 252670 179286
rect 253330 179284 253336 179286
rect 253400 179346 253406 179348
rect 254066 179346 254072 179348
rect 253400 179286 254072 179346
rect 253400 179284 253406 179286
rect 254066 179284 254072 179286
rect 254136 179346 254142 179348
rect 254802 179346 254808 179348
rect 254136 179286 254808 179346
rect 254136 179284 254142 179286
rect 254802 179284 254808 179286
rect 254872 179346 254878 179348
rect 255538 179346 255544 179348
rect 254872 179286 255544 179346
rect 254872 179284 254878 179286
rect 255538 179284 255544 179286
rect 255608 179346 255614 179348
rect 256274 179346 256280 179348
rect 255608 179286 256280 179346
rect 255608 179284 255614 179286
rect 256274 179284 256280 179286
rect 256344 179346 256350 179348
rect 257010 179346 257016 179348
rect 256344 179286 257016 179346
rect 256344 179284 256350 179286
rect 257010 179284 257016 179286
rect 257080 179346 257086 179348
rect 257746 179346 257752 179348
rect 257080 179286 257752 179346
rect 257080 179284 257086 179286
rect 257746 179284 257752 179286
rect 257816 179346 257822 179348
rect 258482 179346 258488 179348
rect 257816 179286 258488 179346
rect 257816 179284 257822 179286
rect 258482 179284 258488 179286
rect 258552 179346 258558 179348
rect 259218 179346 259224 179348
rect 258552 179286 259224 179346
rect 258552 179284 258558 179286
rect 259218 179284 259224 179286
rect 259288 179346 259294 179348
rect 259954 179346 259960 179348
rect 259288 179286 259960 179346
rect 259288 179284 259294 179286
rect 259954 179284 259960 179286
rect 260024 179346 260030 179348
rect 260690 179346 260696 179348
rect 260024 179286 260696 179346
rect 260024 179284 260030 179286
rect 260690 179284 260696 179286
rect 260760 179346 260766 179348
rect 261426 179346 261432 179348
rect 260760 179286 261432 179346
rect 260760 179284 260766 179286
rect 261426 179284 261432 179286
rect 261496 179346 261502 179348
rect 262162 179346 262168 179348
rect 261496 179286 262168 179346
rect 261496 179284 261502 179286
rect 262162 179284 262168 179286
rect 262232 179346 262238 179348
rect 262898 179346 262904 179348
rect 262232 179286 262904 179346
rect 262232 179284 262238 179286
rect 262898 179284 262904 179286
rect 262968 179346 262974 179348
rect 263634 179346 263640 179348
rect 262968 179286 263640 179346
rect 262968 179284 262974 179286
rect 263634 179284 263640 179286
rect 263704 179346 263710 179348
rect 264370 179346 264376 179348
rect 263704 179286 264376 179346
rect 263704 179284 263710 179286
rect 264370 179284 264376 179286
rect 264440 179346 264446 179348
rect 265106 179346 265112 179348
rect 264440 179286 265112 179346
rect 264440 179284 264446 179286
rect 265106 179284 265112 179286
rect 265176 179346 265182 179348
rect 265842 179346 265848 179348
rect 265176 179286 265848 179346
rect 265176 179284 265182 179286
rect 265842 179284 265848 179286
rect 265912 179346 265918 179348
rect 266578 179346 266584 179348
rect 265912 179286 266584 179346
rect 265912 179284 265918 179286
rect 266578 179284 266584 179286
rect 266648 179284 266654 179348
rect 281901 179346 281967 179349
rect 302325 179346 302391 179349
rect 281901 179344 302391 179346
rect 281901 179288 281906 179344
rect 281962 179288 302330 179344
rect 302386 179288 302391 179344
rect 281901 179286 302391 179288
rect 281901 179283 281967 179286
rect 302325 179283 302391 179286
rect 185802 179148 185808 179212
rect 185872 179148 185878 179212
rect 190954 179148 190960 179212
rect 191024 179148 191030 179212
rect 278998 179148 279004 179212
rect 279068 179210 279074 179212
rect 284518 179210 284524 179212
rect 279068 179150 284524 179210
rect 279068 179148 279074 179150
rect 284518 179148 284524 179150
rect 284588 179148 284594 179212
rect 285673 179210 285739 179213
rect 286726 179210 286732 179212
rect 285673 179208 286732 179210
rect 285673 179152 285678 179208
rect 285734 179152 286732 179208
rect 285673 179150 286732 179152
rect 285673 179147 285739 179150
rect 286726 179148 286732 179150
rect 286796 179210 286802 179212
rect 301078 179210 301084 179212
rect 286796 179150 301084 179210
rect 286796 179148 286802 179150
rect 301078 179148 301084 179150
rect 301148 179148 301154 179212
rect 302601 179210 302667 179213
rect 303102 179210 303108 179212
rect 302601 179208 303108 179210
rect 302601 179152 302606 179208
rect 302662 179152 303108 179208
rect 302601 179150 303108 179152
rect 302601 179147 302667 179150
rect 303102 179148 303108 179150
rect 303172 179148 303178 179212
rect 580901 179210 580967 179213
rect 583520 179210 584960 179300
rect 580901 179208 584960 179210
rect 580901 179152 580906 179208
rect 580962 179152 584960 179208
rect 580901 179150 584960 179152
rect 580901 179147 580967 179150
rect 281758 179012 281764 179076
rect 281828 179074 281834 179076
rect 282821 179074 282887 179077
rect 281828 179072 282887 179074
rect 281828 179016 282826 179072
rect 282882 179016 282887 179072
rect 281828 179014 282887 179016
rect 281828 179012 281834 179014
rect 282821 179011 282887 179014
rect 291694 179012 291700 179076
rect 291764 179074 291770 179076
rect 301630 179074 301636 179076
rect 291764 179014 301636 179074
rect 291764 179012 291770 179014
rect 301630 179012 301636 179014
rect 301700 179012 301706 179076
rect 583520 179060 584960 179150
rect 281022 178876 281028 178940
rect 281092 178938 281098 178940
rect 284886 178938 284892 178940
rect 281092 178878 284892 178938
rect 281092 178876 281098 178878
rect 284886 178876 284892 178878
rect 284956 178938 284962 178940
rect 284956 178878 287070 178938
rect 284956 178876 284962 178878
rect 287010 178666 287070 178878
rect 296294 178876 296300 178940
rect 296364 178938 296370 178940
rect 299790 178938 299796 178940
rect 296364 178878 299796 178938
rect 296364 178876 296370 178878
rect 299790 178876 299796 178878
rect 299860 178876 299866 178940
rect 302325 178938 302391 178941
rect 335118 178938 335124 178940
rect 302325 178936 335124 178938
rect 302325 178880 302330 178936
rect 302386 178880 335124 178936
rect 302325 178878 335124 178880
rect 302325 178875 302391 178878
rect 335118 178876 335124 178878
rect 335188 178876 335194 178940
rect 298870 178666 298876 178668
rect 287010 178606 298876 178666
rect 298870 178604 298876 178606
rect 298940 178604 298946 178668
rect 280286 178196 280292 178260
rect 280356 178258 280362 178260
rect 285622 178258 285628 178260
rect 280356 178198 285628 178258
rect 280356 178196 280362 178198
rect 285622 178196 285628 178198
rect 285692 178196 285698 178260
rect 291694 178060 291700 178124
rect 291764 178122 291770 178124
rect 292246 178122 292252 178124
rect 291764 178062 292252 178122
rect 291764 178060 291770 178062
rect 292246 178060 292252 178062
rect 292316 178060 292322 178124
rect 289629 177578 289695 177581
rect 301630 177578 301636 177580
rect 289629 177576 301636 177578
rect 289629 177520 289634 177576
rect 289690 177520 301636 177576
rect 289629 177518 301636 177520
rect 289629 177515 289695 177518
rect 301630 177516 301636 177518
rect 301700 177516 301706 177580
rect 284201 177442 284267 177445
rect 298318 177442 298324 177444
rect 284201 177440 298324 177442
rect 284201 177384 284206 177440
rect 284262 177384 298324 177440
rect 284201 177382 298324 177384
rect 284201 177379 284267 177382
rect 298318 177380 298324 177382
rect 298388 177380 298394 177444
rect 281390 177244 281396 177308
rect 281460 177306 281466 177308
rect 282126 177306 282132 177308
rect 281460 177246 282132 177306
rect 281460 177244 281466 177246
rect 282126 177244 282132 177246
rect 282196 177306 282202 177308
rect 302182 177306 302188 177308
rect 282196 177246 302188 177306
rect 282196 177244 282202 177246
rect 302182 177244 302188 177246
rect 302252 177244 302258 177308
rect 282678 176700 282684 176764
rect 282748 176762 282754 176764
rect 284702 176762 284708 176764
rect 282748 176702 284708 176762
rect 282748 176700 282754 176702
rect 284702 176700 284708 176702
rect 284772 176700 284778 176764
rect 281206 176564 281212 176628
rect 281276 176626 281282 176628
rect 281625 176626 281691 176629
rect 281276 176624 281691 176626
rect 281276 176568 281630 176624
rect 281686 176568 281691 176624
rect 281276 176566 281691 176568
rect 281276 176564 281282 176566
rect 281625 176563 281691 176566
rect 296621 176628 296687 176629
rect 296621 176624 296668 176628
rect 296732 176626 296738 176628
rect 296621 176568 296626 176624
rect 296621 176564 296668 176568
rect 296732 176566 296778 176626
rect 296732 176564 296738 176566
rect 296621 176563 296687 176564
rect -960 175796 480 176036
rect 279550 175340 279556 175404
rect 279620 175402 279626 175404
rect 281942 175402 281948 175404
rect 279620 175342 281948 175402
rect 279620 175340 279626 175342
rect 281942 175340 281948 175342
rect 282012 175340 282018 175404
rect 281942 175204 281948 175268
rect 282012 175266 282018 175268
rect 282862 175266 282868 175268
rect 282012 175206 282868 175266
rect 282012 175204 282018 175206
rect 282862 175204 282868 175206
rect 282932 175204 282938 175268
rect 281441 175130 281507 175133
rect 283557 175130 283623 175133
rect 281441 175128 283623 175130
rect 281441 175072 281446 175128
rect 281502 175072 283562 175128
rect 283618 175072 283623 175128
rect 281441 175070 283623 175072
rect 281441 175067 281507 175070
rect 283557 175067 283623 175070
rect 291142 174524 291148 174588
rect 291212 174586 291218 174588
rect 301814 174586 301820 174588
rect 291212 174526 301820 174586
rect 291212 174524 291218 174526
rect 301814 174524 301820 174526
rect 301884 174524 301890 174588
rect 296621 167108 296687 167109
rect 296621 167106 296668 167108
rect 296576 167104 296668 167106
rect 296576 167048 296626 167104
rect 296576 167046 296668 167048
rect 296621 167044 296668 167046
rect 296732 167044 296738 167108
rect 296621 167043 296687 167044
rect 583520 165732 584960 165972
rect -960 162890 480 162980
rect 3734 162890 3740 162892
rect -960 162830 3740 162890
rect -960 162740 480 162830
rect 3734 162828 3740 162830
rect 3804 162828 3810 162892
rect 296621 161532 296687 161533
rect 296621 161530 296668 161532
rect 296576 161528 296668 161530
rect 296732 161530 296738 161532
rect 296576 161472 296626 161528
rect 296576 161470 296668 161472
rect 296621 161468 296668 161470
rect 296732 161470 296774 161530
rect 296732 161468 296738 161470
rect 296621 161467 296687 161468
rect 296621 161394 296687 161397
rect 296576 161392 296730 161394
rect 296576 161336 296626 161392
rect 296682 161336 296730 161392
rect 296576 161334 296730 161336
rect 296621 161331 296730 161334
rect 296670 161260 296730 161331
rect 296662 161196 296668 161260
rect 296732 161196 296738 161260
rect 281390 157932 281396 157996
rect 281460 157994 281466 157996
rect 304942 157994 304948 157996
rect 281460 157934 304948 157994
rect 281460 157932 281466 157934
rect 304942 157932 304948 157934
rect 305012 157932 305018 157996
rect 301630 157796 301636 157860
rect 301700 157858 301706 157860
rect 311893 157858 311959 157861
rect 301700 157856 311959 157858
rect 301700 157800 311898 157856
rect 311954 157800 311959 157856
rect 301700 157798 311959 157800
rect 301700 157796 301706 157798
rect 311893 157795 311959 157798
rect 284886 157388 284892 157452
rect 284956 157450 284962 157452
rect 286358 157450 286364 157452
rect 284956 157390 286364 157450
rect 284956 157388 284962 157390
rect 286358 157388 286364 157390
rect 286428 157388 286434 157452
rect 303102 157252 303108 157316
rect 303172 157314 303178 157316
rect 306373 157314 306439 157317
rect 303172 157312 306439 157314
rect 303172 157256 306378 157312
rect 306434 157256 306439 157312
rect 303172 157254 306439 157256
rect 303172 157252 303178 157254
rect 306373 157251 306439 157254
rect 300710 156980 300716 157044
rect 300780 157042 300786 157044
rect 309133 157042 309199 157045
rect 300780 157040 309199 157042
rect 300780 156984 309138 157040
rect 309194 156984 309199 157040
rect 300780 156982 309199 156984
rect 300780 156980 300786 156982
rect 309133 156979 309199 156982
rect 296478 156844 296484 156908
rect 296548 156906 296554 156908
rect 306046 156906 306052 156908
rect 296548 156846 306052 156906
rect 296548 156844 296554 156846
rect 306046 156844 306052 156846
rect 306116 156844 306122 156908
rect 292481 156770 292547 156773
rect 304390 156770 304396 156772
rect 292481 156768 304396 156770
rect 292481 156712 292486 156768
rect 292542 156712 304396 156768
rect 292481 156710 304396 156712
rect 292481 156707 292547 156710
rect 304390 156708 304396 156710
rect 304460 156708 304466 156772
rect 284150 156572 284156 156636
rect 284220 156634 284226 156636
rect 300710 156634 300716 156636
rect 284220 156574 300716 156634
rect 284220 156572 284226 156574
rect 300710 156572 300716 156574
rect 300780 156572 300786 156636
rect 301497 156634 301563 156637
rect 303613 156634 303679 156637
rect 301497 156632 303679 156634
rect 301497 156576 301502 156632
rect 301558 156576 303618 156632
rect 303674 156576 303679 156632
rect 301497 156574 303679 156576
rect 301497 156571 301563 156574
rect 303613 156571 303679 156574
rect 304942 156572 304948 156636
rect 305012 156634 305018 156636
rect 314694 156634 314700 156636
rect 305012 156574 314700 156634
rect 305012 156572 305018 156574
rect 314694 156572 314700 156574
rect 314764 156572 314770 156636
rect 301814 155484 301820 155548
rect 301884 155546 301890 155548
rect 313222 155546 313228 155548
rect 301884 155486 313228 155546
rect 301884 155484 301890 155486
rect 313222 155484 313228 155486
rect 313292 155484 313298 155548
rect 284886 155212 284892 155276
rect 284956 155274 284962 155276
rect 335118 155274 335124 155276
rect 284956 155214 335124 155274
rect 284956 155212 284962 155214
rect 335118 155212 335124 155214
rect 335188 155212 335194 155276
rect 300894 153716 300900 153780
rect 300964 153778 300970 153780
rect 315798 153778 315804 153780
rect 300964 153718 315804 153778
rect 300964 153716 300970 153718
rect 315798 153716 315804 153718
rect 315868 153716 315874 153780
rect 580574 152628 580580 152692
rect 580644 152690 580650 152692
rect 583520 152690 584960 152780
rect 580644 152630 584960 152690
rect 580644 152628 580650 152630
rect 583520 152540 584960 152630
rect 296621 151876 296687 151877
rect 296621 151874 296668 151876
rect 296576 151872 296668 151874
rect 296732 151874 296738 151876
rect 296576 151816 296626 151872
rect 296576 151814 296668 151816
rect 296621 151812 296668 151814
rect 296732 151814 296774 151874
rect 296732 151812 296738 151814
rect 296621 151811 296687 151812
rect -960 149834 480 149924
rect 2773 149834 2839 149837
rect -960 149832 2839 149834
rect -960 149776 2778 149832
rect 2834 149776 2839 149832
rect -960 149774 2839 149776
rect -960 149684 480 149774
rect 2773 149771 2839 149774
rect 580574 139300 580580 139364
rect 580644 139362 580650 139364
rect 583520 139362 584960 139452
rect 580644 139302 584960 139362
rect 580644 139300 580650 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 2814 136778 2820 136780
rect -960 136718 2820 136778
rect -960 136628 480 136718
rect 2814 136716 2820 136718
rect 2884 136716 2890 136780
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 580574 112780 580580 112844
rect 580644 112842 580650 112844
rect 583520 112842 584960 112932
rect 580644 112782 584960 112842
rect 580644 112780 580650 112782
rect 583520 112692 584960 112782
rect -960 110516 480 110756
rect 580574 99452 580580 99516
rect 580644 99514 580650 99516
rect 583520 99514 584960 99604
rect 580644 99454 584960 99514
rect 580644 99452 580650 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 2773 97610 2839 97613
rect -960 97608 2839 97610
rect -960 97552 2778 97608
rect 2834 97552 2839 97608
rect -960 97550 2839 97552
rect -960 97460 480 97550
rect 2773 97547 2839 97550
rect 308622 90340 308628 90404
rect 308692 90402 308698 90404
rect 578734 90402 578740 90404
rect 308692 90342 578740 90402
rect 308692 90340 308698 90342
rect 578734 90340 578740 90342
rect 578804 90340 578810 90404
rect 9254 88980 9260 89044
rect 9324 89042 9330 89044
rect 274214 89042 274220 89044
rect 9324 88982 274220 89042
rect 9324 88980 9330 88982
rect 274214 88980 274220 88982
rect 274284 88980 274290 89044
rect 311014 88980 311020 89044
rect 311084 89042 311090 89044
rect 580206 89042 580212 89044
rect 311084 88982 580212 89042
rect 311084 88980 311090 88982
rect 580206 88980 580212 88982
rect 580276 88980 580282 89044
rect 3550 87484 3556 87548
rect 3620 87546 3626 87548
rect 272374 87546 272380 87548
rect 3620 87486 272380 87546
rect 3620 87484 3626 87486
rect 272374 87484 272380 87486
rect 272444 87484 272450 87548
rect 307150 87484 307156 87548
rect 307220 87546 307226 87548
rect 575974 87546 575980 87548
rect 307220 87486 575980 87546
rect 307220 87484 307226 87486
rect 575974 87484 575980 87486
rect 576044 87484 576050 87548
rect 4838 86124 4844 86188
rect 4908 86186 4914 86188
rect 278262 86186 278268 86188
rect 4908 86126 278268 86186
rect 4908 86124 4914 86126
rect 278262 86124 278268 86126
rect 278332 86124 278338 86188
rect 309358 86124 309364 86188
rect 309428 86186 309434 86188
rect 577630 86186 577636 86188
rect 309428 86126 577636 86186
rect 309428 86124 309434 86126
rect 577630 86124 577636 86126
rect 577700 86124 577706 86188
rect 583520 86036 584960 86276
rect -960 84690 480 84780
rect 7598 84764 7604 84828
rect 7668 84826 7674 84828
rect 277158 84826 277164 84828
rect 7668 84766 277164 84826
rect 7668 84764 7674 84766
rect 277158 84764 277164 84766
rect 277228 84764 277234 84828
rect 2773 84690 2839 84693
rect -960 84688 2839 84690
rect -960 84632 2778 84688
rect 2834 84632 2839 84688
rect -960 84630 2839 84632
rect -960 84540 480 84630
rect 2773 84627 2839 84630
rect 6310 83404 6316 83468
rect 6380 83466 6386 83468
rect 276054 83466 276060 83468
rect 6380 83406 276060 83466
rect 6380 83404 6386 83406
rect 276054 83404 276060 83406
rect 276124 83404 276130 83468
rect 6126 82044 6132 82108
rect 6196 82106 6202 82108
rect 276790 82106 276796 82108
rect 6196 82046 276796 82106
rect 6196 82044 6202 82046
rect 276790 82044 276796 82046
rect 276860 82044 276866 82108
rect 7414 80684 7420 80748
rect 7484 80746 7490 80748
rect 277894 80746 277900 80748
rect 7484 80686 277900 80746
rect 7484 80684 7490 80686
rect 277894 80684 277900 80686
rect 277964 80684 277970 80748
rect 6494 77828 6500 77892
rect 6564 77890 6570 77892
rect 274950 77890 274956 77892
rect 6564 77830 274956 77890
rect 6564 77828 6570 77830
rect 274950 77828 274956 77830
rect 275020 77828 275026 77892
rect 3734 76468 3740 76532
rect 3804 76530 3810 76532
rect 273846 76530 273852 76532
rect 3804 76470 273852 76530
rect 3804 76468 3810 76470
rect 273846 76468 273852 76470
rect 273916 76468 273922 76532
rect 7782 75108 7788 75172
rect 7852 75170 7858 75172
rect 275318 75170 275324 75172
rect 7852 75110 275324 75170
rect 7852 75108 7858 75110
rect 275318 75108 275324 75110
rect 275388 75108 275394 75172
rect 308990 75108 308996 75172
rect 309060 75170 309066 75172
rect 577446 75170 577452 75172
rect 309060 75110 577452 75170
rect 309060 75108 309066 75110
rect 577446 75108 577452 75110
rect 577516 75108 577522 75172
rect 9070 73748 9076 73812
rect 9140 73810 9146 73812
rect 276422 73810 276428 73812
rect 9140 73750 276428 73810
rect 9140 73748 9146 73750
rect 276422 73748 276428 73750
rect 276492 73748 276498 73812
rect 580574 72932 580580 72996
rect 580644 72994 580650 72996
rect 583520 72994 584960 73084
rect 580644 72934 584960 72994
rect 580644 72932 580650 72934
rect 583520 72844 584960 72934
rect 4654 72388 4660 72452
rect 4724 72450 4730 72452
rect 277526 72450 277532 72452
rect 4724 72390 277532 72450
rect 4724 72388 4730 72390
rect 277526 72388 277532 72390
rect 277596 72388 277602 72452
rect 307518 72388 307524 72452
rect 307588 72450 307594 72452
rect 576158 72450 576164 72452
rect 307588 72390 576164 72450
rect 307588 72388 307594 72390
rect 576158 72388 576164 72390
rect 576228 72388 576234 72452
rect -960 71634 480 71724
rect 3550 71634 3556 71636
rect -960 71574 3556 71634
rect -960 71484 480 71574
rect 3550 71572 3556 71574
rect 3620 71572 3626 71636
rect 282821 71362 282887 71365
rect 304993 71362 305059 71365
rect 282821 71360 305059 71362
rect 282821 71304 282826 71360
rect 282882 71304 304998 71360
rect 305054 71304 305059 71360
rect 282821 71302 305059 71304
rect 282821 71299 282887 71302
rect 304993 71299 305059 71302
rect 283782 71164 283788 71228
rect 283852 71226 283858 71228
rect 315798 71226 315804 71228
rect 283852 71166 315804 71226
rect 283852 71164 283858 71166
rect 315798 71164 315804 71166
rect 315868 71164 315874 71228
rect 130561 71090 130627 71093
rect 295977 71090 296043 71093
rect 299790 71090 299796 71092
rect 130561 71088 299796 71090
rect 130561 71032 130566 71088
rect 130622 71032 295982 71088
rect 296038 71032 299796 71088
rect 130561 71030 299796 71032
rect 130561 71027 130627 71030
rect 295977 71027 296043 71030
rect 299790 71028 299796 71030
rect 299860 71028 299866 71092
rect 307886 71028 307892 71092
rect 307956 71090 307962 71092
rect 574686 71090 574692 71092
rect 307956 71030 574692 71090
rect 307956 71028 307962 71030
rect 574686 71028 574692 71030
rect 574756 71028 574762 71092
rect 284702 69668 284708 69732
rect 284772 69730 284778 69732
rect 285438 69730 285444 69732
rect 284772 69670 285444 69730
rect 284772 69668 284778 69670
rect 285438 69668 285444 69670
rect 285508 69668 285514 69732
rect 314694 69730 314700 69732
rect 287010 69670 314700 69730
rect 8886 69532 8892 69596
rect 8956 69594 8962 69596
rect 279734 69594 279740 69596
rect 8956 69534 279740 69594
rect 8956 69532 8962 69534
rect 279734 69532 279740 69534
rect 279804 69532 279810 69596
rect 284150 69532 284156 69596
rect 284220 69594 284226 69596
rect 287010 69594 287070 69670
rect 314694 69668 314700 69670
rect 314764 69668 314770 69732
rect 284220 69534 287070 69594
rect 284220 69532 284226 69534
rect 290406 69532 290412 69596
rect 290476 69594 290482 69596
rect 303470 69594 303476 69596
rect 290476 69534 303476 69594
rect 290476 69532 290482 69534
rect 303470 69532 303476 69534
rect 303540 69532 303546 69596
rect 308254 69532 308260 69596
rect 308324 69594 308330 69596
rect 574870 69594 574876 69596
rect 308324 69534 574876 69594
rect 308324 69532 308330 69534
rect 574870 69532 574876 69534
rect 574940 69532 574946 69596
rect 134149 69186 134215 69189
rect 301078 69186 301084 69188
rect 134149 69184 301084 69186
rect 134149 69128 134154 69184
rect 134210 69128 301084 69184
rect 134149 69126 301084 69128
rect 134149 69123 134215 69126
rect 301078 69124 301084 69126
rect 301148 69124 301154 69188
rect 126973 69050 127039 69053
rect 301630 69050 301636 69052
rect 126973 69048 301636 69050
rect 126973 68992 126978 69048
rect 127034 68992 301636 69048
rect 126973 68990 301636 68992
rect 126973 68987 127039 68990
rect 301630 68988 301636 68990
rect 301700 68988 301706 69052
rect 300158 68852 300164 68916
rect 300228 68914 300234 68916
rect 304206 68914 304212 68916
rect 300228 68854 304212 68914
rect 300228 68852 300234 68854
rect 304206 68852 304212 68854
rect 304276 68852 304282 68916
rect 304390 68852 304396 68916
rect 304460 68914 304466 68916
rect 305678 68914 305684 68916
rect 304460 68854 305684 68914
rect 304460 68852 304466 68854
rect 305678 68852 305684 68854
rect 305748 68852 305754 68916
rect 306414 68852 306420 68916
rect 306484 68914 306490 68916
rect 311893 68914 311959 68917
rect 306484 68912 311959 68914
rect 306484 68856 311898 68912
rect 311954 68856 311959 68912
rect 306484 68854 311959 68856
rect 306484 68852 306490 68854
rect 311893 68851 311959 68854
rect 283414 68716 283420 68780
rect 283484 68778 283490 68780
rect 284109 68778 284175 68781
rect 283484 68776 284175 68778
rect 283484 68720 284114 68776
rect 284170 68720 284175 68776
rect 283484 68718 284175 68720
rect 283484 68716 283490 68718
rect 284109 68715 284175 68718
rect 301078 68716 301084 68780
rect 301148 68778 301154 68780
rect 302141 68778 302207 68781
rect 301148 68776 302207 68778
rect 301148 68720 302146 68776
rect 302202 68720 302207 68776
rect 301148 68718 302207 68720
rect 301148 68716 301154 68718
rect 302141 68715 302207 68718
rect 300342 68580 300348 68644
rect 300412 68642 300418 68644
rect 306373 68642 306439 68645
rect 300412 68640 306439 68642
rect 300412 68584 306378 68640
rect 306434 68584 306439 68640
rect 300412 68582 306439 68584
rect 300412 68580 300418 68582
rect 306373 68579 306439 68582
rect 300526 68444 300532 68508
rect 300596 68506 300602 68508
rect 303613 68506 303679 68509
rect 300596 68504 303679 68506
rect 300596 68448 303618 68504
rect 303674 68448 303679 68504
rect 300596 68446 303679 68448
rect 300596 68444 300602 68446
rect 303613 68443 303679 68446
rect 2630 68308 2636 68372
rect 2700 68370 2706 68372
rect 275686 68370 275692 68372
rect 2700 68310 275692 68370
rect 2700 68308 2706 68310
rect 275686 68308 275692 68310
rect 275756 68308 275762 68372
rect 290457 68370 290523 68373
rect 305310 68370 305316 68372
rect 290457 68368 305316 68370
rect 290457 68312 290462 68368
rect 290518 68312 305316 68368
rect 290457 68310 305316 68312
rect 290457 68307 290523 68310
rect 305310 68308 305316 68310
rect 305380 68308 305386 68372
rect 1158 68172 1164 68236
rect 1228 68234 1234 68236
rect 274582 68234 274588 68236
rect 1228 68174 274588 68234
rect 1228 68172 1234 68174
rect 274582 68172 274588 68174
rect 274652 68172 274658 68236
rect 279550 68172 279556 68236
rect 279620 68234 279626 68236
rect 304574 68234 304580 68236
rect 279620 68174 304580 68234
rect 279620 68172 279626 68174
rect 304574 68172 304580 68174
rect 304644 68172 304650 68236
rect 306782 68172 306788 68236
rect 306852 68234 306858 68236
rect 582373 68234 582439 68237
rect 306852 68232 582439 68234
rect 306852 68176 582378 68232
rect 582434 68176 582439 68232
rect 306852 68174 582439 68176
rect 306852 68172 306858 68174
rect 582373 68171 582439 68174
rect 273897 67962 273963 67965
rect 299974 67962 299980 67964
rect 273897 67960 299980 67962
rect 273897 67904 273902 67960
rect 273958 67904 299980 67960
rect 273897 67902 299980 67904
rect 273897 67899 273963 67902
rect 299974 67900 299980 67902
rect 300044 67900 300050 67964
rect 271137 67826 271203 67829
rect 300342 67826 300348 67828
rect 271137 67824 300348 67826
rect 271137 67768 271142 67824
rect 271198 67768 300348 67824
rect 271137 67766 300348 67768
rect 271137 67763 271203 67766
rect 300342 67764 300348 67766
rect 300412 67764 300418 67828
rect 151813 67690 151879 67693
rect 298093 67690 298159 67693
rect 299238 67690 299244 67692
rect 151813 67688 299244 67690
rect 151813 67632 151818 67688
rect 151874 67632 298098 67688
rect 298154 67632 299244 67688
rect 151813 67630 299244 67632
rect 151813 67627 151879 67630
rect 298093 67627 298159 67630
rect 299238 67628 299244 67630
rect 299308 67628 299314 67692
rect 297030 67492 297036 67556
rect 297100 67554 297106 67556
rect 297541 67554 297607 67557
rect 304993 67556 305059 67557
rect 297100 67552 297607 67554
rect 297100 67496 297546 67552
rect 297602 67496 297607 67552
rect 297100 67494 297607 67496
rect 297100 67492 297106 67494
rect 297541 67491 297607 67494
rect 298318 67492 298324 67556
rect 298388 67554 298394 67556
rect 298870 67554 298876 67556
rect 298388 67494 298876 67554
rect 298388 67492 298394 67494
rect 298870 67492 298876 67494
rect 298940 67492 298946 67556
rect 299790 67492 299796 67556
rect 299860 67554 299866 67556
rect 301446 67554 301452 67556
rect 299860 67494 301452 67554
rect 299860 67492 299866 67494
rect 301446 67492 301452 67494
rect 301516 67492 301522 67556
rect 302734 67492 302740 67556
rect 302804 67554 302810 67556
rect 303838 67554 303844 67556
rect 302804 67494 303844 67554
rect 302804 67492 302810 67494
rect 303838 67492 303844 67494
rect 303908 67492 303914 67556
rect 304942 67554 304948 67556
rect 304902 67494 304948 67554
rect 305012 67552 305059 67556
rect 305054 67496 305059 67552
rect 304942 67492 304948 67494
rect 305012 67492 305059 67496
rect 304993 67491 305059 67492
rect 1894 66948 1900 67012
rect 1964 67010 1970 67012
rect 278630 67010 278636 67012
rect 1964 66950 278636 67010
rect 1964 66948 1970 66950
rect 278630 66948 278636 66950
rect 278700 66948 278706 67012
rect 299606 66948 299612 67012
rect 299676 67010 299682 67012
rect 309133 67010 309199 67013
rect 299676 67008 309199 67010
rect 299676 66952 309138 67008
rect 309194 66952 309199 67008
rect 299676 66950 309199 66952
rect 299676 66948 299682 66950
rect 309133 66947 309199 66950
rect 54 66812 60 66876
rect 124 66874 130 66876
rect 279366 66874 279372 66876
rect 124 66814 279372 66874
rect 124 66812 130 66814
rect 279366 66812 279372 66814
rect 279436 66812 279442 66876
rect 302182 66812 302188 66876
rect 302252 66874 302258 66876
rect 313222 66874 313228 66876
rect 302252 66814 313228 66874
rect 302252 66812 302258 66814
rect 313222 66812 313228 66814
rect 313292 66812 313298 66876
rect 279877 66602 279943 66605
rect 299606 66602 299612 66604
rect 279877 66600 299612 66602
rect 279877 66544 279882 66600
rect 279938 66544 299612 66600
rect 279877 66542 299612 66544
rect 279877 66539 279943 66542
rect 299606 66540 299612 66542
rect 299676 66540 299682 66604
rect 274030 66404 274036 66468
rect 274100 66466 274106 66468
rect 298870 66466 298876 66468
rect 274100 66406 298876 66466
rect 274100 66404 274106 66406
rect 298870 66404 298876 66406
rect 298940 66404 298946 66468
rect 158897 66330 158963 66333
rect 298686 66330 298692 66332
rect 158897 66328 298692 66330
rect 158897 66272 158902 66328
rect 158958 66272 298692 66328
rect 158897 66270 298692 66272
rect 158897 66267 158963 66270
rect 298686 66268 298692 66270
rect 298756 66268 298762 66332
rect 137645 65922 137711 65925
rect 300526 65922 300532 65924
rect 137645 65920 300532 65922
rect 137645 65864 137650 65920
rect 137706 65864 300532 65920
rect 137645 65862 300532 65864
rect 137645 65859 137711 65862
rect 300526 65860 300532 65862
rect 300596 65860 300602 65924
rect 148317 65786 148383 65789
rect 279877 65786 279943 65789
rect 148317 65784 279943 65786
rect 148317 65728 148322 65784
rect 148378 65728 279882 65784
rect 279938 65728 279943 65784
rect 148317 65726 279943 65728
rect 148317 65723 148383 65726
rect 279877 65723 279943 65726
rect 3366 65452 3372 65516
rect 3436 65514 3442 65516
rect 272558 65514 272564 65516
rect 3436 65454 272564 65514
rect 3436 65452 3442 65454
rect 272558 65452 272564 65454
rect 272628 65452 272634 65516
rect 144729 64290 144795 64293
rect 273897 64290 273963 64293
rect 144729 64288 273963 64290
rect 144729 64232 144734 64288
rect 144790 64232 273902 64288
rect 273958 64232 273963 64288
rect 144729 64230 273963 64232
rect 144729 64227 144795 64230
rect 273897 64227 273963 64230
rect 141233 64154 141299 64157
rect 271137 64154 271203 64157
rect 141233 64152 271203 64154
rect 141233 64096 141238 64152
rect 141294 64096 271142 64152
rect 271198 64096 271203 64152
rect 141233 64094 271203 64096
rect 141233 64091 141299 64094
rect 271137 64091 271203 64094
rect 155401 62794 155467 62797
rect 274030 62794 274036 62796
rect 155401 62792 274036 62794
rect 155401 62736 155406 62792
rect 155462 62736 274036 62792
rect 155401 62734 274036 62736
rect 155401 62731 155467 62734
rect 274030 62732 274036 62734
rect 274100 62732 274106 62796
rect 580574 59604 580580 59668
rect 580644 59666 580650 59668
rect 583520 59666 584960 59756
rect 580644 59606 584960 59666
rect 580644 59604 580650 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 2773 58578 2839 58581
rect -960 58576 2839 58578
rect -960 58520 2778 58576
rect 2834 58520 2839 58576
rect -960 58518 2839 58520
rect -960 58428 480 58518
rect 2773 58515 2839 58518
rect 583520 46188 584960 46428
rect -960 45522 480 45612
rect 2814 45522 2820 45524
rect -960 45462 2820 45522
rect -960 45372 480 45462
rect 2814 45460 2820 45462
rect 2884 45460 2890 45524
rect 2814 44780 2820 44844
rect 2884 44842 2890 44844
rect 273897 44842 273963 44845
rect 2884 44840 273963 44842
rect 2884 44784 273902 44840
rect 273958 44784 273963 44840
rect 2884 44782 273963 44784
rect 2884 44780 2890 44782
rect 273897 44779 273963 44782
rect 580574 33084 580580 33148
rect 580644 33146 580650 33148
rect 583520 33146 584960 33236
rect 580644 33086 584960 33146
rect 580644 33084 580650 33086
rect 583520 32996 584960 33086
rect -960 32316 480 32556
rect 3550 22612 3556 22676
rect 3620 22674 3626 22676
rect 273294 22674 273300 22676
rect 3620 22614 273300 22674
rect 3620 22612 3626 22614
rect 273294 22612 273300 22614
rect 273364 22612 273370 22676
rect 273897 21994 273963 21997
rect 277710 21994 277716 21996
rect 273897 21992 277716 21994
rect 273897 21936 273902 21992
rect 273958 21936 277716 21992
rect 273897 21934 277716 21936
rect 273897 21931 273963 21934
rect 277710 21932 277716 21934
rect 277780 21994 277786 21996
rect 278681 21994 278747 21997
rect 277780 21992 278747 21994
rect 277780 21936 278686 21992
rect 278742 21936 278747 21992
rect 277780 21934 278747 21936
rect 277780 21932 277786 21934
rect 278681 21931 278747 21934
rect 306414 21932 306420 21996
rect 306484 21994 306490 21996
rect 578918 21994 578924 21996
rect 306484 21934 578924 21994
rect 306484 21932 306490 21934
rect 578918 21932 578924 21934
rect 578988 21932 578994 21996
rect 9438 21796 9444 21860
rect 9508 21858 9514 21860
rect 276606 21858 276612 21860
rect 9508 21798 276612 21858
rect 9508 21796 9514 21798
rect 276606 21796 276612 21798
rect 276676 21796 276682 21860
rect 2078 21660 2084 21724
rect 2148 21722 2154 21724
rect 276238 21722 276244 21724
rect 2148 21662 276244 21722
rect 2148 21660 2154 21662
rect 276238 21660 276244 21662
rect 276308 21660 276314 21724
rect 272558 20572 272564 20636
rect 272628 20634 272634 20636
rect 275686 20634 275692 20636
rect 272628 20574 275692 20634
rect 272628 20572 272634 20574
rect 275686 20572 275692 20574
rect 275756 20572 275762 20636
rect 306598 20572 306604 20636
rect 306668 20634 306674 20636
rect 311014 20634 311020 20636
rect 306668 20574 311020 20634
rect 306668 20572 306674 20574
rect 311014 20572 311020 20574
rect 311084 20572 311090 20636
rect 9857 20498 9923 20501
rect 275318 20498 275324 20500
rect 9857 20496 275324 20498
rect 9857 20440 9862 20496
rect 9918 20440 275324 20496
rect 9857 20438 275324 20440
rect 9857 20435 9923 20438
rect 275318 20436 275324 20438
rect 275388 20436 275394 20500
rect 278681 20498 278747 20501
rect 580574 20498 580580 20500
rect 278681 20496 580580 20498
rect 278681 20440 278686 20496
rect 278742 20440 580580 20496
rect 278681 20438 580580 20440
rect 278681 20435 278747 20438
rect 580574 20436 580580 20438
rect 580644 20498 580650 20500
rect 580644 20438 583586 20498
rect 580644 20436 580650 20438
rect 238 20300 244 20364
rect 308 20362 314 20364
rect 277158 20362 277164 20364
rect 308 20302 277164 20362
rect 308 20300 314 20302
rect 277158 20300 277164 20302
rect 277228 20300 277234 20364
rect 273294 20164 273300 20228
rect 273364 20226 273370 20228
rect 278262 20226 278268 20228
rect 273364 20166 278268 20226
rect 273364 20164 273370 20166
rect 278262 20164 278268 20166
rect 278332 20164 278338 20228
rect 583526 19954 583586 20438
rect 583342 19908 583586 19954
rect 583342 19894 584960 19908
rect 583342 19818 583402 19894
rect 583520 19818 584960 19894
rect 583342 19758 584960 19818
rect 583520 19668 584960 19758
rect 277301 19546 277367 19549
rect 278998 19546 279004 19548
rect 277301 19544 279004 19546
rect -960 19410 480 19500
rect 277301 19488 277306 19544
rect 277362 19488 279004 19544
rect 277301 19486 279004 19488
rect 277301 19483 277367 19486
rect 278998 19484 279004 19486
rect 279068 19484 279074 19548
rect 2773 19410 2839 19413
rect -960 19408 2839 19410
rect -960 19352 2778 19408
rect 2834 19352 2839 19408
rect -960 19350 2839 19352
rect -960 19260 480 19350
rect 2773 19347 2839 19350
rect 277894 19348 277900 19412
rect 277964 19410 277970 19412
rect 278037 19410 278103 19413
rect 277964 19408 278103 19410
rect 277964 19352 278042 19408
rect 278098 19352 278103 19408
rect 277964 19350 278103 19352
rect 277964 19348 277970 19350
rect 278037 19347 278103 19350
rect 273846 19212 273852 19276
rect 273916 19274 273922 19276
rect 278630 19274 278636 19276
rect 273916 19214 278636 19274
rect 273916 19212 273922 19214
rect 278630 19212 278636 19214
rect 278700 19212 278706 19276
rect 272374 19076 272380 19140
rect 272444 19138 272450 19140
rect 277301 19138 277367 19141
rect 272444 19136 277367 19138
rect 272444 19080 277306 19136
rect 277362 19080 277367 19136
rect 272444 19078 277367 19080
rect 272444 19076 272450 19078
rect 277301 19075 277367 19078
rect 5022 18940 5028 19004
rect 5092 19002 5098 19004
rect 276422 19002 276428 19004
rect 5092 18942 276428 19002
rect 5092 18940 5098 18942
rect 276422 18940 276428 18942
rect 276492 18940 276498 19004
rect -960 6490 480 6580
rect 2773 6490 2839 6493
rect -960 6488 2839 6490
rect -960 6432 2778 6488
rect 2834 6432 2839 6488
rect 583520 6476 584960 6716
rect -960 6430 2839 6432
rect -960 6340 480 6430
rect 2773 6427 2839 6430
rect 579797 3498 579863 3501
rect 580758 3498 580764 3500
rect 579797 3496 580764 3498
rect 579797 3440 579802 3496
rect 579858 3440 580764 3496
rect 579797 3438 580764 3440
rect 579797 3435 579863 3438
rect 580758 3436 580764 3438
rect 580828 3436 580834 3500
rect 570321 3362 570387 3365
rect 573909 3362 573975 3365
rect 577405 3362 577471 3365
rect 580901 3362 580967 3365
rect 567150 3360 580967 3362
rect 567150 3304 570326 3360
rect 570382 3304 573914 3360
rect 573970 3304 577410 3360
rect 577466 3304 580906 3360
rect 580962 3304 580967 3360
rect 567150 3302 580967 3304
rect 2773 2818 2839 2821
rect 9949 2818 10015 2821
rect 14733 2818 14799 2821
rect 19425 2818 19491 2821
rect 24209 2818 24275 2821
rect 28901 2818 28967 2821
rect 32397 2818 32463 2821
rect 35985 2818 36051 2821
rect 39573 2818 39639 2821
rect 43069 2818 43135 2821
rect 46657 2818 46723 2821
rect 50153 2818 50219 2821
rect 53741 2818 53807 2821
rect 57237 2818 57303 2821
rect 60825 2818 60891 2821
rect 64321 2818 64387 2821
rect 67909 2818 67975 2821
rect 71497 2818 71563 2821
rect 74993 2818 75059 2821
rect 78581 2818 78647 2821
rect 82077 2818 82143 2821
rect 85665 2818 85731 2821
rect 89161 2818 89227 2821
rect 92749 2818 92815 2821
rect 96245 2818 96311 2821
rect 99833 2818 99899 2821
rect 103329 2818 103395 2821
rect 106917 2818 106983 2821
rect 110505 2818 110571 2821
rect 114001 2818 114067 2821
rect 117589 2818 117655 2821
rect 121085 2818 121151 2821
rect 124673 2818 124739 2821
rect 162485 2818 162551 2821
rect 166073 2818 166139 2821
rect 169569 2818 169635 2821
rect 173157 2818 173223 2821
rect 176653 2818 176719 2821
rect 180241 2818 180307 2821
rect 183737 2818 183803 2821
rect 187325 2818 187391 2821
rect 190821 2818 190887 2821
rect 194409 2818 194475 2821
rect 197905 2818 197971 2821
rect 201493 2818 201559 2821
rect 205081 2818 205147 2821
rect 208577 2818 208643 2821
rect 212165 2818 212231 2821
rect 215661 2818 215727 2821
rect 219249 2818 219315 2821
rect 222745 2818 222811 2821
rect 226333 2818 226399 2821
rect 229829 2818 229895 2821
rect 233417 2818 233483 2821
rect 237005 2818 237071 2821
rect 240501 2818 240567 2821
rect 244089 2818 244155 2821
rect 247585 2818 247651 2821
rect 251173 2818 251239 2821
rect 254669 2818 254735 2821
rect 258257 2818 258323 2821
rect 261753 2818 261819 2821
rect 265341 2818 265407 2821
rect 268837 2818 268903 2821
rect 272425 2818 272491 2821
rect 276013 2818 276079 2821
rect 278037 2818 278103 2821
rect 279509 2818 279575 2821
rect 283097 2818 283163 2821
rect 286593 2818 286659 2821
rect 290181 2818 290247 2821
rect 293677 2818 293743 2821
rect 297265 2818 297331 2821
rect 300761 2818 300827 2821
rect 304349 2818 304415 2821
rect 307937 2818 308003 2821
rect 311433 2818 311499 2821
rect 315021 2818 315087 2821
rect 318517 2818 318583 2821
rect 322105 2818 322171 2821
rect 325601 2818 325667 2821
rect 329189 2818 329255 2821
rect 332685 2818 332751 2821
rect 336273 2818 336339 2821
rect 339861 2818 339927 2821
rect 343357 2818 343423 2821
rect 346945 2818 347011 2821
rect 350441 2818 350507 2821
rect 354029 2818 354095 2821
rect 357525 2818 357591 2821
rect 361113 2818 361179 2821
rect 364609 2818 364675 2821
rect 368197 2818 368263 2821
rect 371693 2818 371759 2821
rect 375281 2818 375347 2821
rect 378869 2818 378935 2821
rect 382365 2818 382431 2821
rect 385953 2818 386019 2821
rect 389449 2818 389515 2821
rect 393037 2818 393103 2821
rect 396533 2818 396599 2821
rect 400121 2818 400187 2821
rect 403617 2818 403683 2821
rect 407205 2818 407271 2821
rect 410793 2818 410859 2821
rect 414289 2818 414355 2821
rect 417877 2818 417943 2821
rect 421373 2818 421439 2821
rect 424961 2818 425027 2821
rect 428457 2818 428523 2821
rect 432045 2818 432111 2821
rect 435541 2818 435607 2821
rect 439129 2818 439195 2821
rect 442625 2818 442691 2821
rect 446213 2818 446279 2821
rect 449801 2818 449867 2821
rect 453297 2818 453363 2821
rect 456885 2818 456951 2821
rect 460381 2818 460447 2821
rect 463969 2818 464035 2821
rect 467465 2818 467531 2821
rect 471053 2818 471119 2821
rect 474549 2818 474615 2821
rect 478137 2818 478203 2821
rect 481725 2818 481791 2821
rect 485221 2818 485287 2821
rect 488809 2818 488875 2821
rect 492305 2818 492371 2821
rect 495893 2818 495959 2821
rect 499389 2818 499455 2821
rect 502977 2818 503043 2821
rect 506473 2818 506539 2821
rect 510061 2818 510127 2821
rect 513557 2818 513623 2821
rect 517145 2818 517211 2821
rect 520733 2818 520799 2821
rect 524229 2818 524295 2821
rect 527817 2818 527883 2821
rect 531313 2818 531379 2821
rect 534901 2818 534967 2821
rect 538397 2818 538463 2821
rect 541985 2818 542051 2821
rect 545481 2818 545547 2821
rect 549069 2818 549135 2821
rect 552657 2818 552723 2821
rect 556153 2818 556219 2821
rect 559741 2818 559807 2821
rect 563237 2818 563303 2821
rect 566825 2818 566891 2821
rect 567150 2818 567210 3302
rect 570321 3299 570387 3302
rect 573909 3299 573975 3302
rect 577405 3299 577471 3302
rect 580901 3299 580967 3302
rect 2773 2816 567210 2818
rect 2773 2760 2778 2816
rect 2834 2760 9954 2816
rect 10010 2760 14738 2816
rect 14794 2760 19430 2816
rect 19486 2760 24214 2816
rect 24270 2760 28906 2816
rect 28962 2760 32402 2816
rect 32458 2760 35990 2816
rect 36046 2760 39578 2816
rect 39634 2760 43074 2816
rect 43130 2760 46662 2816
rect 46718 2760 50158 2816
rect 50214 2760 53746 2816
rect 53802 2760 57242 2816
rect 57298 2760 60830 2816
rect 60886 2760 64326 2816
rect 64382 2760 67914 2816
rect 67970 2760 71502 2816
rect 71558 2760 74998 2816
rect 75054 2760 78586 2816
rect 78642 2760 82082 2816
rect 82138 2760 85670 2816
rect 85726 2760 89166 2816
rect 89222 2760 92754 2816
rect 92810 2760 96250 2816
rect 96306 2760 99838 2816
rect 99894 2760 103334 2816
rect 103390 2760 106922 2816
rect 106978 2760 110510 2816
rect 110566 2760 114006 2816
rect 114062 2760 117594 2816
rect 117650 2760 121090 2816
rect 121146 2760 124678 2816
rect 124734 2760 162490 2816
rect 162546 2760 166078 2816
rect 166134 2760 169574 2816
rect 169630 2760 173162 2816
rect 173218 2760 176658 2816
rect 176714 2760 180246 2816
rect 180302 2760 183742 2816
rect 183798 2760 187330 2816
rect 187386 2760 190826 2816
rect 190882 2760 194414 2816
rect 194470 2760 197910 2816
rect 197966 2760 201498 2816
rect 201554 2760 205086 2816
rect 205142 2760 208582 2816
rect 208638 2760 212170 2816
rect 212226 2760 215666 2816
rect 215722 2760 219254 2816
rect 219310 2760 222750 2816
rect 222806 2760 226338 2816
rect 226394 2760 229834 2816
rect 229890 2760 233422 2816
rect 233478 2760 237010 2816
rect 237066 2760 240506 2816
rect 240562 2760 244094 2816
rect 244150 2760 247590 2816
rect 247646 2760 251178 2816
rect 251234 2760 254674 2816
rect 254730 2760 258262 2816
rect 258318 2760 261758 2816
rect 261814 2760 265346 2816
rect 265402 2760 268842 2816
rect 268898 2760 272430 2816
rect 272486 2760 276018 2816
rect 276074 2760 278042 2816
rect 278098 2760 279514 2816
rect 279570 2760 283102 2816
rect 283158 2760 286598 2816
rect 286654 2760 290186 2816
rect 290242 2760 293682 2816
rect 293738 2760 297270 2816
rect 297326 2760 300766 2816
rect 300822 2760 304354 2816
rect 304410 2760 307942 2816
rect 307998 2760 311438 2816
rect 311494 2760 315026 2816
rect 315082 2760 318522 2816
rect 318578 2760 322110 2816
rect 322166 2760 325606 2816
rect 325662 2760 329194 2816
rect 329250 2760 332690 2816
rect 332746 2760 336278 2816
rect 336334 2760 339866 2816
rect 339922 2760 343362 2816
rect 343418 2760 346950 2816
rect 347006 2760 350446 2816
rect 350502 2760 354034 2816
rect 354090 2760 357530 2816
rect 357586 2760 361118 2816
rect 361174 2760 364614 2816
rect 364670 2760 368202 2816
rect 368258 2760 371698 2816
rect 371754 2760 375286 2816
rect 375342 2760 378874 2816
rect 378930 2760 382370 2816
rect 382426 2760 385958 2816
rect 386014 2760 389454 2816
rect 389510 2760 393042 2816
rect 393098 2760 396538 2816
rect 396594 2760 400126 2816
rect 400182 2760 403622 2816
rect 403678 2760 407210 2816
rect 407266 2760 410798 2816
rect 410854 2760 414294 2816
rect 414350 2760 417882 2816
rect 417938 2760 421378 2816
rect 421434 2760 424966 2816
rect 425022 2760 428462 2816
rect 428518 2760 432050 2816
rect 432106 2760 435546 2816
rect 435602 2760 439134 2816
rect 439190 2760 442630 2816
rect 442686 2760 446218 2816
rect 446274 2760 449806 2816
rect 449862 2760 453302 2816
rect 453358 2760 456890 2816
rect 456946 2760 460386 2816
rect 460442 2760 463974 2816
rect 464030 2760 467470 2816
rect 467526 2760 471058 2816
rect 471114 2760 474554 2816
rect 474610 2760 478142 2816
rect 478198 2760 481730 2816
rect 481786 2760 485226 2816
rect 485282 2760 488814 2816
rect 488870 2760 492310 2816
rect 492366 2760 495898 2816
rect 495954 2760 499394 2816
rect 499450 2760 502982 2816
rect 503038 2760 506478 2816
rect 506534 2760 510066 2816
rect 510122 2760 513562 2816
rect 513618 2760 517150 2816
rect 517206 2760 520738 2816
rect 520794 2760 524234 2816
rect 524290 2760 527822 2816
rect 527878 2760 531318 2816
rect 531374 2760 534906 2816
rect 534962 2760 538402 2816
rect 538458 2760 541990 2816
rect 542046 2760 545486 2816
rect 545542 2760 549074 2816
rect 549130 2760 552662 2816
rect 552718 2760 556158 2816
rect 556214 2760 559746 2816
rect 559802 2760 563242 2816
rect 563298 2760 566830 2816
rect 566886 2760 567210 2816
rect 2773 2758 567210 2760
rect 2773 2755 2839 2758
rect 9949 2755 10015 2758
rect 14733 2755 14799 2758
rect 19425 2755 19491 2758
rect 24209 2755 24275 2758
rect 28901 2755 28967 2758
rect 32397 2755 32463 2758
rect 35985 2755 36051 2758
rect 39573 2755 39639 2758
rect 43069 2755 43135 2758
rect 46657 2755 46723 2758
rect 50153 2755 50219 2758
rect 53741 2755 53807 2758
rect 57237 2755 57303 2758
rect 60825 2755 60891 2758
rect 64321 2755 64387 2758
rect 67909 2755 67975 2758
rect 71497 2755 71563 2758
rect 74993 2755 75059 2758
rect 78581 2755 78647 2758
rect 82077 2755 82143 2758
rect 85665 2755 85731 2758
rect 89161 2755 89227 2758
rect 92749 2755 92815 2758
rect 96245 2755 96311 2758
rect 99833 2755 99899 2758
rect 103329 2755 103395 2758
rect 106917 2755 106983 2758
rect 110505 2755 110571 2758
rect 114001 2755 114067 2758
rect 117589 2755 117655 2758
rect 121085 2755 121151 2758
rect 124673 2755 124739 2758
rect 162485 2755 162551 2758
rect 166073 2755 166139 2758
rect 169569 2755 169635 2758
rect 173157 2755 173223 2758
rect 176653 2755 176719 2758
rect 180241 2755 180307 2758
rect 183737 2755 183803 2758
rect 187325 2755 187391 2758
rect 190821 2755 190887 2758
rect 194409 2755 194475 2758
rect 197905 2755 197971 2758
rect 201493 2755 201559 2758
rect 205081 2755 205147 2758
rect 208577 2755 208643 2758
rect 212165 2755 212231 2758
rect 215661 2755 215727 2758
rect 219249 2755 219315 2758
rect 222745 2755 222811 2758
rect 226333 2755 226399 2758
rect 229829 2755 229895 2758
rect 233417 2755 233483 2758
rect 237005 2755 237071 2758
rect 240501 2755 240567 2758
rect 244089 2755 244155 2758
rect 247585 2755 247651 2758
rect 251173 2755 251239 2758
rect 254669 2755 254735 2758
rect 258257 2755 258323 2758
rect 261753 2755 261819 2758
rect 265341 2755 265407 2758
rect 268837 2755 268903 2758
rect 272425 2755 272491 2758
rect 276013 2755 276079 2758
rect 278037 2755 278103 2758
rect 279509 2755 279575 2758
rect 283097 2755 283163 2758
rect 286593 2755 286659 2758
rect 290181 2755 290247 2758
rect 293677 2755 293743 2758
rect 297265 2755 297331 2758
rect 300761 2755 300827 2758
rect 304349 2755 304415 2758
rect 307937 2755 308003 2758
rect 311433 2755 311499 2758
rect 315021 2755 315087 2758
rect 318517 2755 318583 2758
rect 322105 2755 322171 2758
rect 325601 2755 325667 2758
rect 329189 2755 329255 2758
rect 332685 2755 332751 2758
rect 336273 2755 336339 2758
rect 339861 2755 339927 2758
rect 343357 2755 343423 2758
rect 346945 2755 347011 2758
rect 350441 2755 350507 2758
rect 354029 2755 354095 2758
rect 357525 2755 357591 2758
rect 361113 2755 361179 2758
rect 364609 2755 364675 2758
rect 368197 2755 368263 2758
rect 371693 2755 371759 2758
rect 375281 2755 375347 2758
rect 378869 2755 378935 2758
rect 382365 2755 382431 2758
rect 385953 2755 386019 2758
rect 389449 2755 389515 2758
rect 393037 2755 393103 2758
rect 396533 2755 396599 2758
rect 400121 2755 400187 2758
rect 403617 2755 403683 2758
rect 407205 2755 407271 2758
rect 410793 2755 410859 2758
rect 414289 2755 414355 2758
rect 417877 2755 417943 2758
rect 421373 2755 421439 2758
rect 424961 2755 425027 2758
rect 428457 2755 428523 2758
rect 432045 2755 432111 2758
rect 435541 2755 435607 2758
rect 439129 2755 439195 2758
rect 442625 2755 442691 2758
rect 446213 2755 446279 2758
rect 449801 2755 449867 2758
rect 453297 2755 453363 2758
rect 456885 2755 456951 2758
rect 460381 2755 460447 2758
rect 463969 2755 464035 2758
rect 467465 2755 467531 2758
rect 471053 2755 471119 2758
rect 474549 2755 474615 2758
rect 478137 2755 478203 2758
rect 481725 2755 481791 2758
rect 485221 2755 485287 2758
rect 488809 2755 488875 2758
rect 492305 2755 492371 2758
rect 495893 2755 495959 2758
rect 499389 2755 499455 2758
rect 502977 2755 503043 2758
rect 506473 2755 506539 2758
rect 510061 2755 510127 2758
rect 513557 2755 513623 2758
rect 517145 2755 517211 2758
rect 520733 2755 520799 2758
rect 524229 2755 524295 2758
rect 527817 2755 527883 2758
rect 531313 2755 531379 2758
rect 534901 2755 534967 2758
rect 538397 2755 538463 2758
rect 541985 2755 542051 2758
rect 545481 2755 545547 2758
rect 549069 2755 549135 2758
rect 552657 2755 552723 2758
rect 556153 2755 556219 2758
rect 559741 2755 559807 2758
rect 563237 2755 563303 2758
rect 566825 2755 566891 2758
<< via3 >>
rect 296484 700300 296548 700364
rect 8892 684252 8956 684316
rect 285628 671196 285692 671260
rect 575980 670652 576044 670716
rect 290412 658140 290476 658204
rect 1900 632028 1964 632092
rect 281028 619108 281092 619172
rect 576164 617476 576228 617540
rect 60 605780 124 605844
rect 4660 579940 4724 580004
rect 7420 566884 7484 566948
rect 574692 564300 574756 564364
rect 4844 553828 4908 553892
rect 9076 527852 9140 527916
rect 6132 514796 6196 514860
rect 574876 511260 574940 511324
rect 7604 501740 7668 501804
rect 7788 475628 7852 475692
rect 12388 462572 12452 462636
rect 578740 458084 578804 458148
rect 6316 449516 6380 449580
rect 9260 423540 9324 423604
rect 11100 410484 11164 410548
rect 577452 404908 577516 404972
rect 6500 397428 6564 397492
rect 9812 371316 9876 371380
rect 3372 358396 3436 358460
rect 577636 351868 577700 351932
rect 2084 345340 2148 345404
rect 420958 323444 421022 323508
rect 422182 323444 422246 323508
rect 433334 323444 433398 323508
rect 3556 319228 3620 319292
rect 441660 319228 441724 319292
rect 3740 306172 3804 306236
rect 580212 298692 580276 298756
rect 244 292572 308 292636
rect 281948 281012 282012 281076
rect 287100 280876 287164 280940
rect 284340 280740 284404 280804
rect 300532 276796 300596 276860
rect 302004 275910 302068 275974
rect 301820 273668 301884 273732
rect 301636 272716 301700 272780
rect 3556 271764 3620 271828
rect 5028 271764 5092 271828
rect 300716 270948 300780 271012
rect 300164 269860 300228 269924
rect 300348 268092 300412 268156
rect 3556 267140 3620 267204
rect 580580 259388 580644 259452
rect 441660 259252 441724 259316
rect 580580 258844 580644 258908
rect 441660 253540 441724 253604
rect 301452 249868 301516 249932
rect 300532 249732 300596 249796
rect 302372 249732 302436 249796
rect 299980 248236 300044 248300
rect 300532 247964 300596 248028
rect 300164 247012 300228 247076
rect 578924 245516 578988 245580
rect 3740 242796 3804 242860
rect 9444 242796 9508 242860
rect 2820 241028 2884 241092
rect 301452 239940 301516 240004
rect 304764 239940 304828 240004
rect 441660 239940 441724 240004
rect 425854 239804 425918 239868
rect 337332 237900 337396 237964
rect 425836 237900 425900 237964
rect 300348 237356 300412 237420
rect 308260 237356 308324 237420
rect 329420 236812 329484 236876
rect 353340 236812 353404 236876
rect 312492 236676 312556 236740
rect 324268 236676 324332 236740
rect 325372 236676 325436 236740
rect 350764 236676 350828 236740
rect 323532 236540 323596 236604
rect 336964 236540 337028 236604
rect 349660 236540 349724 236604
rect 408356 236540 408420 236604
rect 337884 236132 337948 236196
rect 340460 236132 340524 236196
rect 299980 235996 300044 236060
rect 305684 235996 305748 236060
rect 316540 235996 316604 236060
rect 318564 235996 318628 236060
rect 319484 235996 319548 236060
rect 322980 235996 323044 236060
rect 323164 235996 323228 236060
rect 325556 235996 325620 236060
rect 334572 235996 334636 236060
rect 336228 235996 336292 236060
rect 340276 235996 340340 236060
rect 344140 235996 344204 236060
rect 300716 235860 300780 235924
rect 308996 235860 309060 235924
rect 323716 235588 323780 235652
rect 338620 235588 338684 235652
rect 313412 235452 313476 235516
rect 333836 235452 333900 235516
rect 333100 235316 333164 235380
rect 366036 235316 366100 235380
rect 320772 235180 320836 235244
rect 356836 235180 356900 235244
rect 325004 234092 325068 234156
rect 343220 234092 343284 234156
rect 78444 233956 78508 234020
rect 90036 233956 90100 234020
rect 318564 233956 318628 234020
rect 350028 233956 350092 234020
rect 89300 233820 89364 233884
rect 110460 233820 110524 233884
rect 301636 233820 301700 233884
rect 309364 233820 309428 233884
rect 310836 233820 310900 233884
rect 323164 233820 323228 233884
rect 327396 233820 327460 233884
rect 363460 233820 363524 233884
rect 317460 232732 317524 232796
rect 346348 232732 346412 232796
rect 321876 232596 321940 232660
rect 360516 232596 360580 232660
rect 301820 232460 301884 232524
rect 309732 232460 309796 232524
rect 314884 232460 314948 232524
rect 338252 232460 338316 232524
rect 338620 232460 338684 232524
rect 400996 232460 401060 232524
rect 315620 231372 315684 231436
rect 337884 231372 337948 231436
rect 318196 231236 318260 231300
rect 348924 231236 348988 231300
rect 360700 231236 360764 231300
rect 370820 231236 370884 231300
rect 326660 231100 326724 231164
rect 361068 231100 361132 231164
rect 326476 230420 326540 230484
rect 333284 230420 333348 230484
rect 315804 230012 315868 230076
rect 342116 230012 342180 230076
rect 321140 229876 321204 229940
rect 358308 229876 358372 229940
rect 306052 229740 306116 229804
rect 320588 229740 320652 229804
rect 333652 229740 333716 229804
rect 405596 229740 405660 229804
rect 315252 228516 315316 228580
rect 339540 228516 339604 228580
rect 327580 228380 327644 228444
rect 356100 228380 356164 228444
rect 317828 228244 317892 228308
rect 347820 228244 347884 228308
rect 356652 228244 356716 228308
rect 395844 228244 395908 228308
rect 317092 227156 317156 227220
rect 345428 227156 345492 227220
rect 321324 227020 321388 227084
rect 359596 227020 359660 227084
rect 314516 226884 314580 226948
rect 323532 226884 323596 226948
rect 331996 226884 332060 226948
rect 386092 226884 386156 226948
rect 311940 225932 312004 225996
rect 329052 225932 329116 225996
rect 340092 225932 340156 225996
rect 348556 225932 348620 225996
rect 324820 225796 324884 225860
rect 346164 225796 346228 225860
rect 316724 225660 316788 225724
rect 340276 225660 340340 225724
rect 328500 225524 328564 225588
rect 368612 225524 368676 225588
rect 307156 224980 307220 225044
rect 312492 224980 312556 225044
rect 324084 224436 324148 224500
rect 341012 224436 341076 224500
rect 307892 224300 307956 224364
rect 319668 224300 319732 224364
rect 331444 224300 331508 224364
rect 391060 224300 391124 224364
rect 312492 224164 312556 224228
rect 327948 224164 328012 224228
rect 328316 224164 328380 224228
rect 331260 224164 331324 224228
rect 332364 224164 332428 224228
rect 398420 224164 398484 224228
rect 322612 223212 322676 223276
rect 330892 223212 330956 223276
rect 330524 223076 330588 223140
rect 343588 223076 343652 223140
rect 323348 222940 323412 223004
rect 334572 222940 334636 223004
rect 334756 222940 334820 223004
rect 373580 222940 373644 223004
rect 311020 222804 311084 222868
rect 322244 222804 322308 222868
rect 330340 222804 330404 222868
rect 383516 222804 383580 222868
rect 334572 221852 334636 221916
rect 349660 221852 349724 221916
rect 313780 221716 313844 221780
rect 334940 221716 335004 221780
rect 322244 221580 322308 221644
rect 361804 221580 361868 221644
rect 313044 221444 313108 221508
rect 332732 221444 332796 221508
rect 333284 221444 333348 221508
rect 403572 221444 403636 221508
rect 320036 220356 320100 220420
rect 354444 220356 354508 220420
rect 320404 220220 320468 220284
rect 355916 220220 355980 220284
rect 307524 220084 307588 220148
rect 316540 220084 316604 220148
rect 329236 220084 329300 220148
rect 375972 220084 376036 220148
rect 324268 218996 324332 219060
rect 336044 218996 336108 219060
rect 580764 218996 580828 219060
rect 326660 218860 326724 218924
rect 358676 218860 358740 218924
rect 319668 218724 319732 218788
rect 353708 218724 353772 218788
rect 302004 218588 302068 218652
rect 309916 218588 309980 218652
rect 311204 218588 311268 218652
rect 327028 218588 327092 218652
rect 331076 218588 331140 218652
rect 388484 218588 388548 218652
rect 318932 217500 318996 217564
rect 351316 217500 351380 217564
rect 300532 217364 300596 217428
rect 305132 217364 305196 217428
rect 319300 217364 319364 217428
rect 352420 217364 352484 217428
rect 306788 217228 306852 217292
rect 319484 217228 319548 217292
rect 329604 217228 329668 217292
rect 378548 217228 378612 217292
rect 330708 217092 330772 217156
rect 331996 217092 332060 217156
rect 325924 216684 325988 216748
rect 329420 216684 329484 216748
rect 324452 216140 324516 216204
rect 330524 216140 330588 216204
rect 332916 216140 332980 216204
rect 338620 216140 338684 216204
rect 306420 216004 306484 216068
rect 311020 216004 311084 216068
rect 314148 216004 314212 216068
rect 324268 216004 324332 216068
rect 312676 215868 312740 215932
rect 328316 216004 328380 216068
rect 328684 216004 328748 216068
rect 360700 216004 360764 216068
rect 329972 215868 330036 215932
rect 381124 215868 381188 215932
rect 333100 215732 333164 215796
rect 316356 215188 316420 215252
rect 325004 215188 325068 215252
rect 325188 214780 325252 214844
rect 340092 214780 340156 214844
rect 332180 214644 332244 214708
rect 356652 214644 356716 214708
rect 281764 214508 281828 214572
rect 312308 214508 312372 214572
rect 330156 214508 330220 214572
rect 331812 214508 331876 214572
rect 393636 214508 393700 214572
rect 302372 213964 302436 214028
rect 310284 213964 310348 214028
rect 10180 213828 10244 213892
rect 12388 213828 12452 213892
rect 1164 213148 1228 213212
rect 11100 213148 11164 213212
rect 326476 213148 326540 213212
rect 311480 213012 311544 213076
rect 312492 213012 312556 213076
rect 322888 213012 322952 213076
rect 326200 213012 326264 213076
rect 327580 213012 327644 213076
rect 328776 213012 328840 213076
rect 334756 213012 334820 213076
rect 308536 212876 308600 212940
rect 327672 212936 327736 212940
rect 327672 212880 327722 212936
rect 327722 212880 327736 212936
rect 327672 212876 327736 212880
rect 281028 193156 281092 193220
rect 284524 193156 284588 193220
rect 78444 192612 78508 192676
rect 90036 192612 90100 192676
rect 89300 192476 89364 192540
rect 110460 192476 110524 192540
rect 301084 191796 301148 191860
rect 335124 191796 335188 191860
rect 337332 191796 337396 191860
rect 2636 190980 2700 191044
rect 10180 190980 10244 191044
rect 298692 190708 298756 190772
rect 281396 190572 281460 190636
rect 282868 190436 282932 190500
rect 291700 190436 291764 190500
rect 298692 190436 298756 190500
rect 9628 190300 9692 190364
rect 283788 189620 283852 189684
rect 299796 189620 299860 189684
rect 283052 189484 283116 189548
rect 299980 189348 300044 189412
rect 282500 189212 282564 189276
rect 292804 189212 292868 189276
rect 283972 189076 284036 189140
rect 285812 188668 285876 188732
rect 301268 188668 301332 188732
rect 284156 188532 284220 188596
rect 296852 188532 296916 188596
rect 302740 188940 302804 189004
rect 302740 188804 302804 188868
rect 292988 188260 293052 188324
rect 300900 188260 300964 188324
rect 302740 188260 302804 188324
rect 302464 188124 302528 188188
rect 291148 187988 291212 188052
rect 283420 187852 283484 187916
rect 292620 187852 292684 187916
rect 301084 187852 301148 187916
rect 301452 187852 301516 187916
rect 299244 187580 299308 187644
rect 299980 187444 300044 187508
rect 281396 187308 281460 187372
rect 283788 187172 283852 187236
rect 299796 187172 299860 187236
rect 300164 187172 300228 187236
rect 300716 187036 300780 187100
rect 284340 186764 284404 186828
rect 297956 186764 298020 186828
rect 283604 186628 283668 186692
rect 297404 186628 297468 186692
rect 299428 186628 299492 186692
rect 298140 186492 298204 186556
rect 297956 186356 298020 186420
rect 283604 186220 283668 186284
rect 299428 186220 299492 186284
rect 283972 186084 284036 186148
rect 284156 185948 284220 186012
rect 296852 185948 296916 186012
rect 296300 185812 296364 185876
rect 299796 185812 299860 185876
rect 295932 185676 295996 185740
rect 295564 185540 295628 185604
rect 295196 185404 295260 185468
rect 294828 185268 294892 185332
rect 294460 185132 294524 185196
rect 294092 184996 294156 185060
rect 283420 184860 283484 184924
rect 287100 184860 287164 184924
rect 292620 184860 292684 184924
rect 293724 184860 293788 184924
rect 282500 184724 282564 184788
rect 292804 184724 292868 184788
rect 293356 184724 293420 184788
rect 282132 184588 282196 184652
rect 299980 184588 300044 184652
rect 300900 184588 300964 184652
rect 292620 184452 292684 184516
rect 282684 184316 282748 184380
rect 301636 184316 301700 184380
rect 291516 184044 291580 184108
rect 290228 183908 290292 183972
rect 290596 183772 290660 183836
rect 291884 183832 291948 183836
rect 291884 183776 291898 183832
rect 291898 183776 291948 183832
rect 291884 183772 291948 183776
rect 300532 183772 300596 183836
rect 289492 183636 289556 183700
rect 289676 183500 289740 183564
rect 288940 183364 289004 183428
rect 289308 183228 289372 183292
rect 289676 183228 289740 183292
rect 288204 183092 288268 183156
rect 287836 182956 287900 183020
rect 287468 182820 287532 182884
rect 287100 182684 287164 182748
rect 301084 182548 301148 182612
rect 281028 182412 281092 182476
rect 300900 182412 300964 182476
rect 285996 182276 286060 182340
rect 285812 182140 285876 182204
rect 288572 182200 288636 182204
rect 288572 182144 288622 182200
rect 288622 182144 288636 182200
rect 288572 182140 288636 182144
rect 301268 182140 301332 182204
rect 285260 182004 285324 182068
rect 285444 181732 285508 181796
rect 281580 181596 281644 181660
rect 284156 181460 284220 181524
rect 283052 181324 283116 181388
rect 283052 181188 283116 181252
rect 284708 181052 284772 181116
rect 281396 180916 281460 180980
rect 302188 180916 302252 180980
rect 282684 180780 282748 180844
rect 281580 180644 281644 180708
rect 282132 180372 282196 180436
rect 292988 180372 293052 180436
rect 296852 180372 296916 180436
rect 290596 180236 290660 180300
rect 300532 180236 300596 180300
rect 300164 180100 300228 180164
rect 302556 179828 302620 179892
rect 298876 179692 298940 179756
rect 300900 179692 300964 179756
rect 299244 179556 299308 179620
rect 290044 179420 290108 179484
rect 290596 179420 290660 179484
rect 182128 179284 182192 179348
rect 182864 179284 182928 179348
rect 183600 179284 183664 179348
rect 184336 179284 184400 179348
rect 185072 179284 185136 179348
rect 186544 179284 186608 179348
rect 187280 179284 187344 179348
rect 188016 179284 188080 179348
rect 188752 179284 188816 179348
rect 189488 179284 189552 179348
rect 190224 179284 190288 179348
rect 191696 179284 191760 179348
rect 192432 179284 192496 179348
rect 193168 179284 193232 179348
rect 193904 179284 193968 179348
rect 194640 179284 194704 179348
rect 195376 179284 195440 179348
rect 196112 179284 196176 179348
rect 196848 179284 196912 179348
rect 197584 179284 197648 179348
rect 198320 179284 198384 179348
rect 214788 179284 214852 179348
rect 215524 179284 215588 179348
rect 216260 179284 216324 179348
rect 216996 179284 217060 179348
rect 217732 179284 217796 179348
rect 218468 179284 218532 179348
rect 219204 179284 219268 179348
rect 219940 179284 220004 179348
rect 220860 179284 220924 179348
rect 221412 179284 221476 179348
rect 222148 179284 222212 179348
rect 222884 179284 222948 179348
rect 223620 179284 223684 179348
rect 248920 179284 248984 179348
rect 249656 179284 249720 179348
rect 250392 179284 250456 179348
rect 251128 179284 251192 179348
rect 251864 179284 251928 179348
rect 252600 179284 252664 179348
rect 253336 179284 253400 179348
rect 254072 179284 254136 179348
rect 254808 179284 254872 179348
rect 255544 179284 255608 179348
rect 256280 179284 256344 179348
rect 257016 179284 257080 179348
rect 257752 179284 257816 179348
rect 258488 179284 258552 179348
rect 259224 179284 259288 179348
rect 259960 179284 260024 179348
rect 260696 179284 260760 179348
rect 261432 179284 261496 179348
rect 262168 179284 262232 179348
rect 262904 179284 262968 179348
rect 263640 179284 263704 179348
rect 264376 179284 264440 179348
rect 265112 179284 265176 179348
rect 265848 179284 265912 179348
rect 266584 179284 266648 179348
rect 185808 179148 185872 179212
rect 190960 179148 191024 179212
rect 279004 179148 279068 179212
rect 284524 179148 284588 179212
rect 286732 179148 286796 179212
rect 301084 179148 301148 179212
rect 303108 179148 303172 179212
rect 281764 179012 281828 179076
rect 291700 179012 291764 179076
rect 301636 179012 301700 179076
rect 281028 178876 281092 178940
rect 284892 178876 284956 178940
rect 296300 178876 296364 178940
rect 299796 178876 299860 178940
rect 335124 178876 335188 178940
rect 298876 178604 298940 178668
rect 280292 178196 280356 178260
rect 285628 178196 285692 178260
rect 291700 178060 291764 178124
rect 292252 178060 292316 178124
rect 301636 177516 301700 177580
rect 298324 177380 298388 177444
rect 281396 177244 281460 177308
rect 282132 177244 282196 177308
rect 302188 177244 302252 177308
rect 282684 176700 282748 176764
rect 284708 176700 284772 176764
rect 281212 176564 281276 176628
rect 296668 176624 296732 176628
rect 296668 176568 296682 176624
rect 296682 176568 296732 176624
rect 296668 176564 296732 176568
rect 279556 175340 279620 175404
rect 281948 175340 282012 175404
rect 281948 175204 282012 175268
rect 282868 175204 282932 175268
rect 291148 174524 291212 174588
rect 301820 174524 301884 174588
rect 296668 167104 296732 167108
rect 296668 167048 296682 167104
rect 296682 167048 296732 167104
rect 296668 167044 296732 167048
rect 3740 162828 3804 162892
rect 296668 161528 296732 161532
rect 296668 161472 296682 161528
rect 296682 161472 296732 161528
rect 296668 161468 296732 161472
rect 296668 161196 296732 161260
rect 281396 157932 281460 157996
rect 304948 157932 305012 157996
rect 301636 157796 301700 157860
rect 284892 157388 284956 157452
rect 286364 157388 286428 157452
rect 303108 157252 303172 157316
rect 300716 156980 300780 157044
rect 296484 156844 296548 156908
rect 306052 156844 306116 156908
rect 304396 156708 304460 156772
rect 284156 156572 284220 156636
rect 300716 156572 300780 156636
rect 304948 156572 305012 156636
rect 314700 156572 314764 156636
rect 301820 155484 301884 155548
rect 313228 155484 313292 155548
rect 284892 155212 284956 155276
rect 335124 155212 335188 155276
rect 300900 153716 300964 153780
rect 315804 153716 315868 153780
rect 580580 152628 580644 152692
rect 296668 151872 296732 151876
rect 296668 151816 296682 151872
rect 296682 151816 296732 151872
rect 296668 151812 296732 151816
rect 580580 139300 580644 139364
rect 2820 136716 2884 136780
rect 580580 112780 580644 112844
rect 580580 99452 580644 99516
rect 308628 90340 308692 90404
rect 578740 90340 578804 90404
rect 9260 88980 9324 89044
rect 274220 88980 274284 89044
rect 311020 88980 311084 89044
rect 580212 88980 580276 89044
rect 3556 87484 3620 87548
rect 272380 87484 272444 87548
rect 307156 87484 307220 87548
rect 575980 87484 576044 87548
rect 4844 86124 4908 86188
rect 278268 86124 278332 86188
rect 309364 86124 309428 86188
rect 577636 86124 577700 86188
rect 7604 84764 7668 84828
rect 277164 84764 277228 84828
rect 6316 83404 6380 83468
rect 276060 83404 276124 83468
rect 6132 82044 6196 82108
rect 276796 82044 276860 82108
rect 7420 80684 7484 80748
rect 277900 80684 277964 80748
rect 6500 77828 6564 77892
rect 274956 77828 275020 77892
rect 3740 76468 3804 76532
rect 273852 76468 273916 76532
rect 7788 75108 7852 75172
rect 275324 75108 275388 75172
rect 308996 75108 309060 75172
rect 577452 75108 577516 75172
rect 9076 73748 9140 73812
rect 276428 73748 276492 73812
rect 580580 72932 580644 72996
rect 4660 72388 4724 72452
rect 277532 72388 277596 72452
rect 307524 72388 307588 72452
rect 576164 72388 576228 72452
rect 3556 71572 3620 71636
rect 283788 71164 283852 71228
rect 315804 71164 315868 71228
rect 299796 71028 299860 71092
rect 307892 71028 307956 71092
rect 574692 71028 574756 71092
rect 284708 69668 284772 69732
rect 285444 69668 285508 69732
rect 8892 69532 8956 69596
rect 279740 69532 279804 69596
rect 284156 69532 284220 69596
rect 314700 69668 314764 69732
rect 290412 69532 290476 69596
rect 303476 69532 303540 69596
rect 308260 69532 308324 69596
rect 574876 69532 574940 69596
rect 301084 69124 301148 69188
rect 301636 68988 301700 69052
rect 300164 68852 300228 68916
rect 304212 68852 304276 68916
rect 304396 68852 304460 68916
rect 305684 68852 305748 68916
rect 306420 68852 306484 68916
rect 283420 68716 283484 68780
rect 301084 68716 301148 68780
rect 300348 68580 300412 68644
rect 300532 68444 300596 68508
rect 2636 68308 2700 68372
rect 275692 68308 275756 68372
rect 305316 68308 305380 68372
rect 1164 68172 1228 68236
rect 274588 68172 274652 68236
rect 279556 68172 279620 68236
rect 304580 68172 304644 68236
rect 306788 68172 306852 68236
rect 299980 67900 300044 67964
rect 300348 67764 300412 67828
rect 299244 67628 299308 67692
rect 297036 67492 297100 67556
rect 298324 67492 298388 67556
rect 298876 67492 298940 67556
rect 299796 67492 299860 67556
rect 301452 67492 301516 67556
rect 302740 67492 302804 67556
rect 303844 67492 303908 67556
rect 304948 67552 305012 67556
rect 304948 67496 304998 67552
rect 304998 67496 305012 67552
rect 304948 67492 305012 67496
rect 1900 66948 1964 67012
rect 278636 66948 278700 67012
rect 299612 66948 299676 67012
rect 60 66812 124 66876
rect 279372 66812 279436 66876
rect 302188 66812 302252 66876
rect 313228 66812 313292 66876
rect 299612 66540 299676 66604
rect 274036 66404 274100 66468
rect 298876 66404 298940 66468
rect 298692 66268 298756 66332
rect 300532 65860 300596 65924
rect 3372 65452 3436 65516
rect 272564 65452 272628 65516
rect 274036 62732 274100 62796
rect 580580 59604 580644 59668
rect 2820 45460 2884 45524
rect 2820 44780 2884 44844
rect 580580 33084 580644 33148
rect 3556 22612 3620 22676
rect 273300 22612 273364 22676
rect 277716 21932 277780 21996
rect 306420 21932 306484 21996
rect 578924 21932 578988 21996
rect 9444 21796 9508 21860
rect 276612 21796 276676 21860
rect 2084 21660 2148 21724
rect 276244 21660 276308 21724
rect 272564 20572 272628 20636
rect 275692 20572 275756 20636
rect 306604 20572 306668 20636
rect 311020 20572 311084 20636
rect 275324 20436 275388 20500
rect 580580 20436 580644 20500
rect 244 20300 308 20364
rect 277164 20300 277228 20364
rect 273300 20164 273364 20228
rect 278268 20164 278332 20228
rect 279004 19484 279068 19548
rect 277900 19348 277964 19412
rect 273852 19212 273916 19276
rect 278636 19212 278700 19276
rect 272380 19076 272444 19140
rect 5028 18940 5092 19004
rect 276428 18940 276492 19004
rect 580764 3436 580828 3500
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 -7066 -8106 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 -6106 -7146 710042
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 -5146 -6186 709082
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 -4186 -5226 708122
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 -3226 -4266 707162
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 -2266 -3306 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 694454 -2346 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 694218 -2934 694454
rect -2698 694218 -2614 694454
rect -2378 694218 -2346 694454
rect -2966 694134 -2346 694218
rect -2966 693898 -2934 694134
rect -2698 693898 -2614 694134
rect -2378 693898 -2346 694134
rect -2966 684454 -2346 693898
rect -2966 684218 -2934 684454
rect -2698 684218 -2614 684454
rect -2378 684218 -2346 684454
rect -2966 684134 -2346 684218
rect -2966 683898 -2934 684134
rect -2698 683898 -2614 684134
rect -2378 683898 -2346 684134
rect -2966 674454 -2346 683898
rect -2966 674218 -2934 674454
rect -2698 674218 -2614 674454
rect -2378 674218 -2346 674454
rect -2966 674134 -2346 674218
rect -2966 673898 -2934 674134
rect -2698 673898 -2614 674134
rect -2378 673898 -2346 674134
rect -2966 664454 -2346 673898
rect -2966 664218 -2934 664454
rect -2698 664218 -2614 664454
rect -2378 664218 -2346 664454
rect -2966 664134 -2346 664218
rect -2966 663898 -2934 664134
rect -2698 663898 -2614 664134
rect -2378 663898 -2346 664134
rect -2966 654454 -2346 663898
rect -2966 654218 -2934 654454
rect -2698 654218 -2614 654454
rect -2378 654218 -2346 654454
rect -2966 654134 -2346 654218
rect -2966 653898 -2934 654134
rect -2698 653898 -2614 654134
rect -2378 653898 -2346 654134
rect -2966 644454 -2346 653898
rect -2966 644218 -2934 644454
rect -2698 644218 -2614 644454
rect -2378 644218 -2346 644454
rect -2966 644134 -2346 644218
rect -2966 643898 -2934 644134
rect -2698 643898 -2614 644134
rect -2378 643898 -2346 644134
rect -2966 634454 -2346 643898
rect -2966 634218 -2934 634454
rect -2698 634218 -2614 634454
rect -2378 634218 -2346 634454
rect -2966 634134 -2346 634218
rect -2966 633898 -2934 634134
rect -2698 633898 -2614 634134
rect -2378 633898 -2346 634134
rect -2966 624454 -2346 633898
rect -2966 624218 -2934 624454
rect -2698 624218 -2614 624454
rect -2378 624218 -2346 624454
rect -2966 624134 -2346 624218
rect -2966 623898 -2934 624134
rect -2698 623898 -2614 624134
rect -2378 623898 -2346 624134
rect -2966 614454 -2346 623898
rect -2966 614218 -2934 614454
rect -2698 614218 -2614 614454
rect -2378 614218 -2346 614454
rect -2966 614134 -2346 614218
rect -2966 613898 -2934 614134
rect -2698 613898 -2614 614134
rect -2378 613898 -2346 614134
rect -2966 604454 -2346 613898
rect -2966 604218 -2934 604454
rect -2698 604218 -2614 604454
rect -2378 604218 -2346 604454
rect -2966 604134 -2346 604218
rect -2966 603898 -2934 604134
rect -2698 603898 -2614 604134
rect -2378 603898 -2346 604134
rect -2966 594454 -2346 603898
rect -2966 594218 -2934 594454
rect -2698 594218 -2614 594454
rect -2378 594218 -2346 594454
rect -2966 594134 -2346 594218
rect -2966 593898 -2934 594134
rect -2698 593898 -2614 594134
rect -2378 593898 -2346 594134
rect -2966 584454 -2346 593898
rect -2966 584218 -2934 584454
rect -2698 584218 -2614 584454
rect -2378 584218 -2346 584454
rect -2966 584134 -2346 584218
rect -2966 583898 -2934 584134
rect -2698 583898 -2614 584134
rect -2378 583898 -2346 584134
rect -2966 574454 -2346 583898
rect -2966 574218 -2934 574454
rect -2698 574218 -2614 574454
rect -2378 574218 -2346 574454
rect -2966 574134 -2346 574218
rect -2966 573898 -2934 574134
rect -2698 573898 -2614 574134
rect -2378 573898 -2346 574134
rect -2966 564454 -2346 573898
rect -2966 564218 -2934 564454
rect -2698 564218 -2614 564454
rect -2378 564218 -2346 564454
rect -2966 564134 -2346 564218
rect -2966 563898 -2934 564134
rect -2698 563898 -2614 564134
rect -2378 563898 -2346 564134
rect -2966 554454 -2346 563898
rect -2966 554218 -2934 554454
rect -2698 554218 -2614 554454
rect -2378 554218 -2346 554454
rect -2966 554134 -2346 554218
rect -2966 553898 -2934 554134
rect -2698 553898 -2614 554134
rect -2378 553898 -2346 554134
rect -2966 544454 -2346 553898
rect -2966 544218 -2934 544454
rect -2698 544218 -2614 544454
rect -2378 544218 -2346 544454
rect -2966 544134 -2346 544218
rect -2966 543898 -2934 544134
rect -2698 543898 -2614 544134
rect -2378 543898 -2346 544134
rect -2966 534454 -2346 543898
rect -2966 534218 -2934 534454
rect -2698 534218 -2614 534454
rect -2378 534218 -2346 534454
rect -2966 534134 -2346 534218
rect -2966 533898 -2934 534134
rect -2698 533898 -2614 534134
rect -2378 533898 -2346 534134
rect -2966 524454 -2346 533898
rect -2966 524218 -2934 524454
rect -2698 524218 -2614 524454
rect -2378 524218 -2346 524454
rect -2966 524134 -2346 524218
rect -2966 523898 -2934 524134
rect -2698 523898 -2614 524134
rect -2378 523898 -2346 524134
rect -2966 514454 -2346 523898
rect -2966 514218 -2934 514454
rect -2698 514218 -2614 514454
rect -2378 514218 -2346 514454
rect -2966 514134 -2346 514218
rect -2966 513898 -2934 514134
rect -2698 513898 -2614 514134
rect -2378 513898 -2346 514134
rect -2966 504454 -2346 513898
rect -2966 504218 -2934 504454
rect -2698 504218 -2614 504454
rect -2378 504218 -2346 504454
rect -2966 504134 -2346 504218
rect -2966 503898 -2934 504134
rect -2698 503898 -2614 504134
rect -2378 503898 -2346 504134
rect -2966 494454 -2346 503898
rect -2966 494218 -2934 494454
rect -2698 494218 -2614 494454
rect -2378 494218 -2346 494454
rect -2966 494134 -2346 494218
rect -2966 493898 -2934 494134
rect -2698 493898 -2614 494134
rect -2378 493898 -2346 494134
rect -2966 484454 -2346 493898
rect -2966 484218 -2934 484454
rect -2698 484218 -2614 484454
rect -2378 484218 -2346 484454
rect -2966 484134 -2346 484218
rect -2966 483898 -2934 484134
rect -2698 483898 -2614 484134
rect -2378 483898 -2346 484134
rect -2966 474454 -2346 483898
rect -2966 474218 -2934 474454
rect -2698 474218 -2614 474454
rect -2378 474218 -2346 474454
rect -2966 474134 -2346 474218
rect -2966 473898 -2934 474134
rect -2698 473898 -2614 474134
rect -2378 473898 -2346 474134
rect -2966 464454 -2346 473898
rect -2966 464218 -2934 464454
rect -2698 464218 -2614 464454
rect -2378 464218 -2346 464454
rect -2966 464134 -2346 464218
rect -2966 463898 -2934 464134
rect -2698 463898 -2614 464134
rect -2378 463898 -2346 464134
rect -2966 454454 -2346 463898
rect -2966 454218 -2934 454454
rect -2698 454218 -2614 454454
rect -2378 454218 -2346 454454
rect -2966 454134 -2346 454218
rect -2966 453898 -2934 454134
rect -2698 453898 -2614 454134
rect -2378 453898 -2346 454134
rect -2966 444454 -2346 453898
rect -2966 444218 -2934 444454
rect -2698 444218 -2614 444454
rect -2378 444218 -2346 444454
rect -2966 444134 -2346 444218
rect -2966 443898 -2934 444134
rect -2698 443898 -2614 444134
rect -2378 443898 -2346 444134
rect -2966 434454 -2346 443898
rect -2966 434218 -2934 434454
rect -2698 434218 -2614 434454
rect -2378 434218 -2346 434454
rect -2966 434134 -2346 434218
rect -2966 433898 -2934 434134
rect -2698 433898 -2614 434134
rect -2378 433898 -2346 434134
rect -2966 424454 -2346 433898
rect -2966 424218 -2934 424454
rect -2698 424218 -2614 424454
rect -2378 424218 -2346 424454
rect -2966 424134 -2346 424218
rect -2966 423898 -2934 424134
rect -2698 423898 -2614 424134
rect -2378 423898 -2346 424134
rect -2966 414454 -2346 423898
rect -2966 414218 -2934 414454
rect -2698 414218 -2614 414454
rect -2378 414218 -2346 414454
rect -2966 414134 -2346 414218
rect -2966 413898 -2934 414134
rect -2698 413898 -2614 414134
rect -2378 413898 -2346 414134
rect -2966 404454 -2346 413898
rect -2966 404218 -2934 404454
rect -2698 404218 -2614 404454
rect -2378 404218 -2346 404454
rect -2966 404134 -2346 404218
rect -2966 403898 -2934 404134
rect -2698 403898 -2614 404134
rect -2378 403898 -2346 404134
rect -2966 394454 -2346 403898
rect -2966 394218 -2934 394454
rect -2698 394218 -2614 394454
rect -2378 394218 -2346 394454
rect -2966 394134 -2346 394218
rect -2966 393898 -2934 394134
rect -2698 393898 -2614 394134
rect -2378 393898 -2346 394134
rect -2966 384454 -2346 393898
rect -2966 384218 -2934 384454
rect -2698 384218 -2614 384454
rect -2378 384218 -2346 384454
rect -2966 384134 -2346 384218
rect -2966 383898 -2934 384134
rect -2698 383898 -2614 384134
rect -2378 383898 -2346 384134
rect -2966 374454 -2346 383898
rect -2966 374218 -2934 374454
rect -2698 374218 -2614 374454
rect -2378 374218 -2346 374454
rect -2966 374134 -2346 374218
rect -2966 373898 -2934 374134
rect -2698 373898 -2614 374134
rect -2378 373898 -2346 374134
rect -2966 364454 -2346 373898
rect -2966 364218 -2934 364454
rect -2698 364218 -2614 364454
rect -2378 364218 -2346 364454
rect -2966 364134 -2346 364218
rect -2966 363898 -2934 364134
rect -2698 363898 -2614 364134
rect -2378 363898 -2346 364134
rect -2966 354454 -2346 363898
rect -2966 354218 -2934 354454
rect -2698 354218 -2614 354454
rect -2378 354218 -2346 354454
rect -2966 354134 -2346 354218
rect -2966 353898 -2934 354134
rect -2698 353898 -2614 354134
rect -2378 353898 -2346 354134
rect -2966 344454 -2346 353898
rect -2966 344218 -2934 344454
rect -2698 344218 -2614 344454
rect -2378 344218 -2346 344454
rect -2966 344134 -2346 344218
rect -2966 343898 -2934 344134
rect -2698 343898 -2614 344134
rect -2378 343898 -2346 344134
rect -2966 334454 -2346 343898
rect -2966 334218 -2934 334454
rect -2698 334218 -2614 334454
rect -2378 334218 -2346 334454
rect -2966 334134 -2346 334218
rect -2966 333898 -2934 334134
rect -2698 333898 -2614 334134
rect -2378 333898 -2346 334134
rect -2966 324454 -2346 333898
rect -2966 324218 -2934 324454
rect -2698 324218 -2614 324454
rect -2378 324218 -2346 324454
rect -2966 324134 -2346 324218
rect -2966 323898 -2934 324134
rect -2698 323898 -2614 324134
rect -2378 323898 -2346 324134
rect -2966 314454 -2346 323898
rect -2966 314218 -2934 314454
rect -2698 314218 -2614 314454
rect -2378 314218 -2346 314454
rect -2966 314134 -2346 314218
rect -2966 313898 -2934 314134
rect -2698 313898 -2614 314134
rect -2378 313898 -2346 314134
rect -2966 304454 -2346 313898
rect -2966 304218 -2934 304454
rect -2698 304218 -2614 304454
rect -2378 304218 -2346 304454
rect -2966 304134 -2346 304218
rect -2966 303898 -2934 304134
rect -2698 303898 -2614 304134
rect -2378 303898 -2346 304134
rect -2966 294454 -2346 303898
rect -2966 294218 -2934 294454
rect -2698 294218 -2614 294454
rect -2378 294218 -2346 294454
rect -2966 294134 -2346 294218
rect -2966 293898 -2934 294134
rect -2698 293898 -2614 294134
rect -2378 293898 -2346 294134
rect -2966 284454 -2346 293898
rect -2966 284218 -2934 284454
rect -2698 284218 -2614 284454
rect -2378 284218 -2346 284454
rect -2966 284134 -2346 284218
rect -2966 283898 -2934 284134
rect -2698 283898 -2614 284134
rect -2378 283898 -2346 284134
rect -2966 274454 -2346 283898
rect -2966 274218 -2934 274454
rect -2698 274218 -2614 274454
rect -2378 274218 -2346 274454
rect -2966 274134 -2346 274218
rect -2966 273898 -2934 274134
rect -2698 273898 -2614 274134
rect -2378 273898 -2346 274134
rect -2966 264454 -2346 273898
rect -2966 264218 -2934 264454
rect -2698 264218 -2614 264454
rect -2378 264218 -2346 264454
rect -2966 264134 -2346 264218
rect -2966 263898 -2934 264134
rect -2698 263898 -2614 264134
rect -2378 263898 -2346 264134
rect -2966 254454 -2346 263898
rect -2966 254218 -2934 254454
rect -2698 254218 -2614 254454
rect -2378 254218 -2346 254454
rect -2966 254134 -2346 254218
rect -2966 253898 -2934 254134
rect -2698 253898 -2614 254134
rect -2378 253898 -2346 254134
rect -2966 244454 -2346 253898
rect -2966 244218 -2934 244454
rect -2698 244218 -2614 244454
rect -2378 244218 -2346 244454
rect -2966 244134 -2346 244218
rect -2966 243898 -2934 244134
rect -2698 243898 -2614 244134
rect -2378 243898 -2346 244134
rect -2966 234454 -2346 243898
rect -2966 234218 -2934 234454
rect -2698 234218 -2614 234454
rect -2378 234218 -2346 234454
rect -2966 234134 -2346 234218
rect -2966 233898 -2934 234134
rect -2698 233898 -2614 234134
rect -2378 233898 -2346 234134
rect -2966 224454 -2346 233898
rect -2966 224218 -2934 224454
rect -2698 224218 -2614 224454
rect -2378 224218 -2346 224454
rect -2966 224134 -2346 224218
rect -2966 223898 -2934 224134
rect -2698 223898 -2614 224134
rect -2378 223898 -2346 224134
rect -2966 214454 -2346 223898
rect -2966 214218 -2934 214454
rect -2698 214218 -2614 214454
rect -2378 214218 -2346 214454
rect -2966 214134 -2346 214218
rect -2966 213898 -2934 214134
rect -2698 213898 -2614 214134
rect -2378 213898 -2346 214134
rect -2966 204454 -2346 213898
rect -2966 204218 -2934 204454
rect -2698 204218 -2614 204454
rect -2378 204218 -2346 204454
rect -2966 204134 -2346 204218
rect -2966 203898 -2934 204134
rect -2698 203898 -2614 204134
rect -2378 203898 -2346 204134
rect -2966 194454 -2346 203898
rect -2966 194218 -2934 194454
rect -2698 194218 -2614 194454
rect -2378 194218 -2346 194454
rect -2966 194134 -2346 194218
rect -2966 193898 -2934 194134
rect -2698 193898 -2614 194134
rect -2378 193898 -2346 194134
rect -2966 184454 -2346 193898
rect -2966 184218 -2934 184454
rect -2698 184218 -2614 184454
rect -2378 184218 -2346 184454
rect -2966 184134 -2346 184218
rect -2966 183898 -2934 184134
rect -2698 183898 -2614 184134
rect -2378 183898 -2346 184134
rect -2966 174454 -2346 183898
rect -2966 174218 -2934 174454
rect -2698 174218 -2614 174454
rect -2378 174218 -2346 174454
rect -2966 174134 -2346 174218
rect -2966 173898 -2934 174134
rect -2698 173898 -2614 174134
rect -2378 173898 -2346 174134
rect -2966 164454 -2346 173898
rect -2966 164218 -2934 164454
rect -2698 164218 -2614 164454
rect -2378 164218 -2346 164454
rect -2966 164134 -2346 164218
rect -2966 163898 -2934 164134
rect -2698 163898 -2614 164134
rect -2378 163898 -2346 164134
rect -2966 154454 -2346 163898
rect -2966 154218 -2934 154454
rect -2698 154218 -2614 154454
rect -2378 154218 -2346 154454
rect -2966 154134 -2346 154218
rect -2966 153898 -2934 154134
rect -2698 153898 -2614 154134
rect -2378 153898 -2346 154134
rect -2966 144454 -2346 153898
rect -2966 144218 -2934 144454
rect -2698 144218 -2614 144454
rect -2378 144218 -2346 144454
rect -2966 144134 -2346 144218
rect -2966 143898 -2934 144134
rect -2698 143898 -2614 144134
rect -2378 143898 -2346 144134
rect -2966 134454 -2346 143898
rect -2966 134218 -2934 134454
rect -2698 134218 -2614 134454
rect -2378 134218 -2346 134454
rect -2966 134134 -2346 134218
rect -2966 133898 -2934 134134
rect -2698 133898 -2614 134134
rect -2378 133898 -2346 134134
rect -2966 124454 -2346 133898
rect -2966 124218 -2934 124454
rect -2698 124218 -2614 124454
rect -2378 124218 -2346 124454
rect -2966 124134 -2346 124218
rect -2966 123898 -2934 124134
rect -2698 123898 -2614 124134
rect -2378 123898 -2346 124134
rect -2966 114454 -2346 123898
rect -2966 114218 -2934 114454
rect -2698 114218 -2614 114454
rect -2378 114218 -2346 114454
rect -2966 114134 -2346 114218
rect -2966 113898 -2934 114134
rect -2698 113898 -2614 114134
rect -2378 113898 -2346 114134
rect -2966 104454 -2346 113898
rect -2966 104218 -2934 104454
rect -2698 104218 -2614 104454
rect -2378 104218 -2346 104454
rect -2966 104134 -2346 104218
rect -2966 103898 -2934 104134
rect -2698 103898 -2614 104134
rect -2378 103898 -2346 104134
rect -2966 94454 -2346 103898
rect -2966 94218 -2934 94454
rect -2698 94218 -2614 94454
rect -2378 94218 -2346 94454
rect -2966 94134 -2346 94218
rect -2966 93898 -2934 94134
rect -2698 93898 -2614 94134
rect -2378 93898 -2346 94134
rect -2966 84454 -2346 93898
rect -2966 84218 -2934 84454
rect -2698 84218 -2614 84454
rect -2378 84218 -2346 84454
rect -2966 84134 -2346 84218
rect -2966 83898 -2934 84134
rect -2698 83898 -2614 84134
rect -2378 83898 -2346 84134
rect -2966 74454 -2346 83898
rect -2966 74218 -2934 74454
rect -2698 74218 -2614 74454
rect -2378 74218 -2346 74454
rect -2966 74134 -2346 74218
rect -2966 73898 -2934 74134
rect -2698 73898 -2614 74134
rect -2378 73898 -2346 74134
rect -2966 64454 -2346 73898
rect -2966 64218 -2934 64454
rect -2698 64218 -2614 64454
rect -2378 64218 -2346 64454
rect -2966 64134 -2346 64218
rect -2966 63898 -2934 64134
rect -2698 63898 -2614 64134
rect -2378 63898 -2346 64134
rect -2966 54454 -2346 63898
rect -2966 54218 -2934 54454
rect -2698 54218 -2614 54454
rect -2378 54218 -2346 54454
rect -2966 54134 -2346 54218
rect -2966 53898 -2934 54134
rect -2698 53898 -2614 54134
rect -2378 53898 -2346 54134
rect -2966 44454 -2346 53898
rect -2966 44218 -2934 44454
rect -2698 44218 -2614 44454
rect -2378 44218 -2346 44454
rect -2966 44134 -2346 44218
rect -2966 43898 -2934 44134
rect -2698 43898 -2614 44134
rect -2378 43898 -2346 44134
rect -2966 34454 -2346 43898
rect -2966 34218 -2934 34454
rect -2698 34218 -2614 34454
rect -2378 34218 -2346 34454
rect -2966 34134 -2346 34218
rect -2966 33898 -2934 34134
rect -2698 33898 -2614 34134
rect -2378 33898 -2346 34134
rect -2966 -1306 -2346 33898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 698174 -1386 704282
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 296483 700364 296549 700365
rect 296483 700300 296484 700364
rect 296548 700300 296549 700364
rect 296483 700299 296549 700300
rect -2006 697938 -1974 698174
rect -1738 697938 -1654 698174
rect -1418 697938 -1386 698174
rect -2006 697854 -1386 697938
rect -2006 697618 -1974 697854
rect -1738 697618 -1654 697854
rect -1418 697618 -1386 697854
rect -2006 688174 -1386 697618
rect -2006 687938 -1974 688174
rect -1738 687938 -1654 688174
rect -1418 687938 -1386 688174
rect -2006 687854 -1386 687938
rect -2006 687618 -1974 687854
rect -1738 687618 -1654 687854
rect -1418 687618 -1386 687854
rect -2006 678174 -1386 687618
rect 8891 684316 8957 684317
rect 8891 684252 8892 684316
rect 8956 684252 8957 684316
rect 8891 684251 8957 684252
rect -2006 677938 -1974 678174
rect -1738 677938 -1654 678174
rect -1418 677938 -1386 678174
rect -2006 677854 -1386 677938
rect -2006 677618 -1974 677854
rect -1738 677618 -1654 677854
rect -1418 677618 -1386 677854
rect -2006 668174 -1386 677618
rect -2006 667938 -1974 668174
rect -1738 667938 -1654 668174
rect -1418 667938 -1386 668174
rect -2006 667854 -1386 667938
rect -2006 667618 -1974 667854
rect -1738 667618 -1654 667854
rect -1418 667618 -1386 667854
rect -2006 658174 -1386 667618
rect -2006 657938 -1974 658174
rect -1738 657938 -1654 658174
rect -1418 657938 -1386 658174
rect -2006 657854 -1386 657938
rect -2006 657618 -1974 657854
rect -1738 657618 -1654 657854
rect -1418 657618 -1386 657854
rect -2006 648174 -1386 657618
rect -2006 647938 -1974 648174
rect -1738 647938 -1654 648174
rect -1418 647938 -1386 648174
rect -2006 647854 -1386 647938
rect -2006 647618 -1974 647854
rect -1738 647618 -1654 647854
rect -1418 647618 -1386 647854
rect -2006 638174 -1386 647618
rect -2006 637938 -1974 638174
rect -1738 637938 -1654 638174
rect -1418 637938 -1386 638174
rect -2006 637854 -1386 637938
rect -2006 637618 -1974 637854
rect -1738 637618 -1654 637854
rect -1418 637618 -1386 637854
rect -2006 628174 -1386 637618
rect 1899 632092 1965 632093
rect 1899 632028 1900 632092
rect 1964 632028 1965 632092
rect 1899 632027 1965 632028
rect -2006 627938 -1974 628174
rect -1738 627938 -1654 628174
rect -1418 627938 -1386 628174
rect -2006 627854 -1386 627938
rect -2006 627618 -1974 627854
rect -1738 627618 -1654 627854
rect -1418 627618 -1386 627854
rect -2006 618174 -1386 627618
rect -2006 617938 -1974 618174
rect -1738 617938 -1654 618174
rect -1418 617938 -1386 618174
rect -2006 617854 -1386 617938
rect -2006 617618 -1974 617854
rect -1738 617618 -1654 617854
rect -1418 617618 -1386 617854
rect -2006 608174 -1386 617618
rect -2006 607938 -1974 608174
rect -1738 607938 -1654 608174
rect -1418 607938 -1386 608174
rect -2006 607854 -1386 607938
rect -2006 607618 -1974 607854
rect -1738 607618 -1654 607854
rect -1418 607618 -1386 607854
rect -2006 598174 -1386 607618
rect 59 605844 125 605845
rect 59 605780 60 605844
rect 124 605780 125 605844
rect 59 605779 125 605780
rect -2006 597938 -1974 598174
rect -1738 597938 -1654 598174
rect -1418 597938 -1386 598174
rect -2006 597854 -1386 597938
rect -2006 597618 -1974 597854
rect -1738 597618 -1654 597854
rect -1418 597618 -1386 597854
rect -2006 588174 -1386 597618
rect -2006 587938 -1974 588174
rect -1738 587938 -1654 588174
rect -1418 587938 -1386 588174
rect -2006 587854 -1386 587938
rect -2006 587618 -1974 587854
rect -1738 587618 -1654 587854
rect -1418 587618 -1386 587854
rect -2006 578174 -1386 587618
rect -2006 577938 -1974 578174
rect -1738 577938 -1654 578174
rect -1418 577938 -1386 578174
rect -2006 577854 -1386 577938
rect -2006 577618 -1974 577854
rect -1738 577618 -1654 577854
rect -1418 577618 -1386 577854
rect -2006 568174 -1386 577618
rect -2006 567938 -1974 568174
rect -1738 567938 -1654 568174
rect -1418 567938 -1386 568174
rect -2006 567854 -1386 567938
rect -2006 567618 -1974 567854
rect -1738 567618 -1654 567854
rect -1418 567618 -1386 567854
rect -2006 558174 -1386 567618
rect -2006 557938 -1974 558174
rect -1738 557938 -1654 558174
rect -1418 557938 -1386 558174
rect -2006 557854 -1386 557938
rect -2006 557618 -1974 557854
rect -1738 557618 -1654 557854
rect -1418 557618 -1386 557854
rect -2006 548174 -1386 557618
rect -2006 547938 -1974 548174
rect -1738 547938 -1654 548174
rect -1418 547938 -1386 548174
rect -2006 547854 -1386 547938
rect -2006 547618 -1974 547854
rect -1738 547618 -1654 547854
rect -1418 547618 -1386 547854
rect -2006 538174 -1386 547618
rect -2006 537938 -1974 538174
rect -1738 537938 -1654 538174
rect -1418 537938 -1386 538174
rect -2006 537854 -1386 537938
rect -2006 537618 -1974 537854
rect -1738 537618 -1654 537854
rect -1418 537618 -1386 537854
rect -2006 528174 -1386 537618
rect -2006 527938 -1974 528174
rect -1738 527938 -1654 528174
rect -1418 527938 -1386 528174
rect -2006 527854 -1386 527938
rect -2006 527618 -1974 527854
rect -1738 527618 -1654 527854
rect -1418 527618 -1386 527854
rect -2006 518174 -1386 527618
rect -2006 517938 -1974 518174
rect -1738 517938 -1654 518174
rect -1418 517938 -1386 518174
rect -2006 517854 -1386 517938
rect -2006 517618 -1974 517854
rect -1738 517618 -1654 517854
rect -1418 517618 -1386 517854
rect -2006 508174 -1386 517618
rect -2006 507938 -1974 508174
rect -1738 507938 -1654 508174
rect -1418 507938 -1386 508174
rect -2006 507854 -1386 507938
rect -2006 507618 -1974 507854
rect -1738 507618 -1654 507854
rect -1418 507618 -1386 507854
rect -2006 498174 -1386 507618
rect -2006 497938 -1974 498174
rect -1738 497938 -1654 498174
rect -1418 497938 -1386 498174
rect -2006 497854 -1386 497938
rect -2006 497618 -1974 497854
rect -1738 497618 -1654 497854
rect -1418 497618 -1386 497854
rect -2006 488174 -1386 497618
rect -2006 487938 -1974 488174
rect -1738 487938 -1654 488174
rect -1418 487938 -1386 488174
rect -2006 487854 -1386 487938
rect -2006 487618 -1974 487854
rect -1738 487618 -1654 487854
rect -1418 487618 -1386 487854
rect -2006 478174 -1386 487618
rect -2006 477938 -1974 478174
rect -1738 477938 -1654 478174
rect -1418 477938 -1386 478174
rect -2006 477854 -1386 477938
rect -2006 477618 -1974 477854
rect -1738 477618 -1654 477854
rect -1418 477618 -1386 477854
rect -2006 468174 -1386 477618
rect -2006 467938 -1974 468174
rect -1738 467938 -1654 468174
rect -1418 467938 -1386 468174
rect -2006 467854 -1386 467938
rect -2006 467618 -1974 467854
rect -1738 467618 -1654 467854
rect -1418 467618 -1386 467854
rect -2006 458174 -1386 467618
rect -2006 457938 -1974 458174
rect -1738 457938 -1654 458174
rect -1418 457938 -1386 458174
rect -2006 457854 -1386 457938
rect -2006 457618 -1974 457854
rect -1738 457618 -1654 457854
rect -1418 457618 -1386 457854
rect -2006 448174 -1386 457618
rect -2006 447938 -1974 448174
rect -1738 447938 -1654 448174
rect -1418 447938 -1386 448174
rect -2006 447854 -1386 447938
rect -2006 447618 -1974 447854
rect -1738 447618 -1654 447854
rect -1418 447618 -1386 447854
rect -2006 438174 -1386 447618
rect -2006 437938 -1974 438174
rect -1738 437938 -1654 438174
rect -1418 437938 -1386 438174
rect -2006 437854 -1386 437938
rect -2006 437618 -1974 437854
rect -1738 437618 -1654 437854
rect -1418 437618 -1386 437854
rect -2006 428174 -1386 437618
rect -2006 427938 -1974 428174
rect -1738 427938 -1654 428174
rect -1418 427938 -1386 428174
rect -2006 427854 -1386 427938
rect -2006 427618 -1974 427854
rect -1738 427618 -1654 427854
rect -1418 427618 -1386 427854
rect -2006 418174 -1386 427618
rect -2006 417938 -1974 418174
rect -1738 417938 -1654 418174
rect -1418 417938 -1386 418174
rect -2006 417854 -1386 417938
rect -2006 417618 -1974 417854
rect -1738 417618 -1654 417854
rect -1418 417618 -1386 417854
rect -2006 408174 -1386 417618
rect -2006 407938 -1974 408174
rect -1738 407938 -1654 408174
rect -1418 407938 -1386 408174
rect -2006 407854 -1386 407938
rect -2006 407618 -1974 407854
rect -1738 407618 -1654 407854
rect -1418 407618 -1386 407854
rect -2006 398174 -1386 407618
rect -2006 397938 -1974 398174
rect -1738 397938 -1654 398174
rect -1418 397938 -1386 398174
rect -2006 397854 -1386 397938
rect -2006 397618 -1974 397854
rect -1738 397618 -1654 397854
rect -1418 397618 -1386 397854
rect -2006 388174 -1386 397618
rect -2006 387938 -1974 388174
rect -1738 387938 -1654 388174
rect -1418 387938 -1386 388174
rect -2006 387854 -1386 387938
rect -2006 387618 -1974 387854
rect -1738 387618 -1654 387854
rect -1418 387618 -1386 387854
rect -2006 378174 -1386 387618
rect -2006 377938 -1974 378174
rect -1738 377938 -1654 378174
rect -1418 377938 -1386 378174
rect -2006 377854 -1386 377938
rect -2006 377618 -1974 377854
rect -1738 377618 -1654 377854
rect -1418 377618 -1386 377854
rect -2006 368174 -1386 377618
rect -2006 367938 -1974 368174
rect -1738 367938 -1654 368174
rect -1418 367938 -1386 368174
rect -2006 367854 -1386 367938
rect -2006 367618 -1974 367854
rect -1738 367618 -1654 367854
rect -1418 367618 -1386 367854
rect -2006 358174 -1386 367618
rect -2006 357938 -1974 358174
rect -1738 357938 -1654 358174
rect -1418 357938 -1386 358174
rect -2006 357854 -1386 357938
rect -2006 357618 -1974 357854
rect -1738 357618 -1654 357854
rect -1418 357618 -1386 357854
rect -2006 348174 -1386 357618
rect -2006 347938 -1974 348174
rect -1738 347938 -1654 348174
rect -1418 347938 -1386 348174
rect -2006 347854 -1386 347938
rect -2006 347618 -1974 347854
rect -1738 347618 -1654 347854
rect -1418 347618 -1386 347854
rect -2006 338174 -1386 347618
rect -2006 337938 -1974 338174
rect -1738 337938 -1654 338174
rect -1418 337938 -1386 338174
rect -2006 337854 -1386 337938
rect -2006 337618 -1974 337854
rect -1738 337618 -1654 337854
rect -1418 337618 -1386 337854
rect -2006 328174 -1386 337618
rect -2006 327938 -1974 328174
rect -1738 327938 -1654 328174
rect -1418 327938 -1386 328174
rect -2006 327854 -1386 327938
rect -2006 327618 -1974 327854
rect -1738 327618 -1654 327854
rect -1418 327618 -1386 327854
rect -2006 318174 -1386 327618
rect -2006 317938 -1974 318174
rect -1738 317938 -1654 318174
rect -1418 317938 -1386 318174
rect -2006 317854 -1386 317938
rect -2006 317618 -1974 317854
rect -1738 317618 -1654 317854
rect -1418 317618 -1386 317854
rect -2006 308174 -1386 317618
rect -2006 307938 -1974 308174
rect -1738 307938 -1654 308174
rect -1418 307938 -1386 308174
rect -2006 307854 -1386 307938
rect -2006 307618 -1974 307854
rect -1738 307618 -1654 307854
rect -1418 307618 -1386 307854
rect -2006 298174 -1386 307618
rect -2006 297938 -1974 298174
rect -1738 297938 -1654 298174
rect -1418 297938 -1386 298174
rect -2006 297854 -1386 297938
rect -2006 297618 -1974 297854
rect -1738 297618 -1654 297854
rect -1418 297618 -1386 297854
rect -2006 288174 -1386 297618
rect -2006 287938 -1974 288174
rect -1738 287938 -1654 288174
rect -1418 287938 -1386 288174
rect -2006 287854 -1386 287938
rect -2006 287618 -1974 287854
rect -1738 287618 -1654 287854
rect -1418 287618 -1386 287854
rect -2006 278174 -1386 287618
rect -2006 277938 -1974 278174
rect -1738 277938 -1654 278174
rect -1418 277938 -1386 278174
rect -2006 277854 -1386 277938
rect -2006 277618 -1974 277854
rect -1738 277618 -1654 277854
rect -1418 277618 -1386 277854
rect -2006 268174 -1386 277618
rect -2006 267938 -1974 268174
rect -1738 267938 -1654 268174
rect -1418 267938 -1386 268174
rect -2006 267854 -1386 267938
rect -2006 267618 -1974 267854
rect -1738 267618 -1654 267854
rect -1418 267618 -1386 267854
rect -2006 258174 -1386 267618
rect -2006 257938 -1974 258174
rect -1738 257938 -1654 258174
rect -1418 257938 -1386 258174
rect -2006 257854 -1386 257938
rect -2006 257618 -1974 257854
rect -1738 257618 -1654 257854
rect -1418 257618 -1386 257854
rect -2006 248174 -1386 257618
rect -2006 247938 -1974 248174
rect -1738 247938 -1654 248174
rect -1418 247938 -1386 248174
rect -2006 247854 -1386 247938
rect -2006 247618 -1974 247854
rect -1738 247618 -1654 247854
rect -1418 247618 -1386 247854
rect -2006 238174 -1386 247618
rect -2006 237938 -1974 238174
rect -1738 237938 -1654 238174
rect -1418 237938 -1386 238174
rect -2006 237854 -1386 237938
rect -2006 237618 -1974 237854
rect -1738 237618 -1654 237854
rect -1418 237618 -1386 237854
rect -2006 228174 -1386 237618
rect -2006 227938 -1974 228174
rect -1738 227938 -1654 228174
rect -1418 227938 -1386 228174
rect -2006 227854 -1386 227938
rect -2006 227618 -1974 227854
rect -1738 227618 -1654 227854
rect -1418 227618 -1386 227854
rect -2006 218174 -1386 227618
rect -2006 217938 -1974 218174
rect -1738 217938 -1654 218174
rect -1418 217938 -1386 218174
rect -2006 217854 -1386 217938
rect -2006 217618 -1974 217854
rect -1738 217618 -1654 217854
rect -1418 217618 -1386 217854
rect -2006 208174 -1386 217618
rect -2006 207938 -1974 208174
rect -1738 207938 -1654 208174
rect -1418 207938 -1386 208174
rect -2006 207854 -1386 207938
rect -2006 207618 -1974 207854
rect -1738 207618 -1654 207854
rect -1418 207618 -1386 207854
rect -2006 198174 -1386 207618
rect -2006 197938 -1974 198174
rect -1738 197938 -1654 198174
rect -1418 197938 -1386 198174
rect -2006 197854 -1386 197938
rect -2006 197618 -1974 197854
rect -1738 197618 -1654 197854
rect -1418 197618 -1386 197854
rect -2006 188174 -1386 197618
rect -2006 187938 -1974 188174
rect -1738 187938 -1654 188174
rect -1418 187938 -1386 188174
rect -2006 187854 -1386 187938
rect -2006 187618 -1974 187854
rect -1738 187618 -1654 187854
rect -1418 187618 -1386 187854
rect -2006 178174 -1386 187618
rect -2006 177938 -1974 178174
rect -1738 177938 -1654 178174
rect -1418 177938 -1386 178174
rect -2006 177854 -1386 177938
rect -2006 177618 -1974 177854
rect -1738 177618 -1654 177854
rect -1418 177618 -1386 177854
rect -2006 168174 -1386 177618
rect -2006 167938 -1974 168174
rect -1738 167938 -1654 168174
rect -1418 167938 -1386 168174
rect -2006 167854 -1386 167938
rect -2006 167618 -1974 167854
rect -1738 167618 -1654 167854
rect -1418 167618 -1386 167854
rect -2006 158174 -1386 167618
rect -2006 157938 -1974 158174
rect -1738 157938 -1654 158174
rect -1418 157938 -1386 158174
rect -2006 157854 -1386 157938
rect -2006 157618 -1974 157854
rect -1738 157618 -1654 157854
rect -1418 157618 -1386 157854
rect -2006 148174 -1386 157618
rect -2006 147938 -1974 148174
rect -1738 147938 -1654 148174
rect -1418 147938 -1386 148174
rect -2006 147854 -1386 147938
rect -2006 147618 -1974 147854
rect -1738 147618 -1654 147854
rect -1418 147618 -1386 147854
rect -2006 138174 -1386 147618
rect -2006 137938 -1974 138174
rect -1738 137938 -1654 138174
rect -1418 137938 -1386 138174
rect -2006 137854 -1386 137938
rect -2006 137618 -1974 137854
rect -1738 137618 -1654 137854
rect -1418 137618 -1386 137854
rect -2006 128174 -1386 137618
rect -2006 127938 -1974 128174
rect -1738 127938 -1654 128174
rect -1418 127938 -1386 128174
rect -2006 127854 -1386 127938
rect -2006 127618 -1974 127854
rect -1738 127618 -1654 127854
rect -1418 127618 -1386 127854
rect -2006 118174 -1386 127618
rect -2006 117938 -1974 118174
rect -1738 117938 -1654 118174
rect -1418 117938 -1386 118174
rect -2006 117854 -1386 117938
rect -2006 117618 -1974 117854
rect -1738 117618 -1654 117854
rect -1418 117618 -1386 117854
rect -2006 108174 -1386 117618
rect -2006 107938 -1974 108174
rect -1738 107938 -1654 108174
rect -1418 107938 -1386 108174
rect -2006 107854 -1386 107938
rect -2006 107618 -1974 107854
rect -1738 107618 -1654 107854
rect -1418 107618 -1386 107854
rect -2006 98174 -1386 107618
rect -2006 97938 -1974 98174
rect -1738 97938 -1654 98174
rect -1418 97938 -1386 98174
rect -2006 97854 -1386 97938
rect -2006 97618 -1974 97854
rect -1738 97618 -1654 97854
rect -1418 97618 -1386 97854
rect -2006 88174 -1386 97618
rect -2006 87938 -1974 88174
rect -1738 87938 -1654 88174
rect -1418 87938 -1386 88174
rect -2006 87854 -1386 87938
rect -2006 87618 -1974 87854
rect -1738 87618 -1654 87854
rect -1418 87618 -1386 87854
rect -2006 78174 -1386 87618
rect -2006 77938 -1974 78174
rect -1738 77938 -1654 78174
rect -1418 77938 -1386 78174
rect -2006 77854 -1386 77938
rect -2006 77618 -1974 77854
rect -1738 77618 -1654 77854
rect -1418 77618 -1386 77854
rect -2006 68174 -1386 77618
rect -2006 67938 -1974 68174
rect -1738 67938 -1654 68174
rect -1418 67938 -1386 68174
rect -2006 67854 -1386 67938
rect -2006 67618 -1974 67854
rect -1738 67618 -1654 67854
rect -1418 67618 -1386 67854
rect -2006 58174 -1386 67618
rect 62 66877 122 605779
rect 243 292636 309 292637
rect 243 292572 244 292636
rect 308 292572 309 292636
rect 243 292571 309 292572
rect 59 66876 125 66877
rect 59 66812 60 66876
rect 124 66812 125 66876
rect 59 66811 125 66812
rect -2006 57938 -1974 58174
rect -1738 57938 -1654 58174
rect -1418 57938 -1386 58174
rect -2006 57854 -1386 57938
rect -2006 57618 -1974 57854
rect -1738 57618 -1654 57854
rect -1418 57618 -1386 57854
rect -2006 48174 -1386 57618
rect -2006 47938 -1974 48174
rect -1738 47938 -1654 48174
rect -1418 47938 -1386 48174
rect -2006 47854 -1386 47938
rect -2006 47618 -1974 47854
rect -1738 47618 -1654 47854
rect -1418 47618 -1386 47854
rect -2006 38174 -1386 47618
rect -2006 37938 -1974 38174
rect -1738 37938 -1654 38174
rect -1418 37938 -1386 38174
rect -2006 37854 -1386 37938
rect -2006 37618 -1974 37854
rect -1738 37618 -1654 37854
rect -1418 37618 -1386 37854
rect -2006 -346 -1386 37618
rect 246 20365 306 292571
rect 1163 213212 1229 213213
rect 1163 213148 1164 213212
rect 1228 213148 1229 213212
rect 1163 213147 1229 213148
rect 1166 68237 1226 213147
rect 1163 68236 1229 68237
rect 1163 68172 1164 68236
rect 1228 68172 1229 68236
rect 1163 68171 1229 68172
rect 1902 67013 1962 632027
rect 4659 580004 4725 580005
rect 4659 579940 4660 580004
rect 4724 579940 4725 580004
rect 4659 579939 4725 579940
rect 3371 358460 3437 358461
rect 3371 358396 3372 358460
rect 3436 358396 3437 358460
rect 3371 358395 3437 358396
rect 2083 345404 2149 345405
rect 2083 345340 2084 345404
rect 2148 345340 2149 345404
rect 2083 345339 2149 345340
rect 1899 67012 1965 67013
rect 1899 66948 1900 67012
rect 1964 66948 1965 67012
rect 1899 66947 1965 66948
rect 2086 21725 2146 345339
rect 2819 241092 2885 241093
rect 2819 241028 2820 241092
rect 2884 241028 2885 241092
rect 2819 241027 2885 241028
rect 2635 191044 2701 191045
rect 2635 190980 2636 191044
rect 2700 190980 2701 191044
rect 2635 190979 2701 190980
rect 2638 68373 2698 190979
rect 2822 136781 2882 241027
rect 2819 136780 2885 136781
rect 2819 136716 2820 136780
rect 2884 136716 2885 136780
rect 2819 136715 2885 136716
rect 2635 68372 2701 68373
rect 2635 68308 2636 68372
rect 2700 68308 2701 68372
rect 2635 68307 2701 68308
rect 2822 45525 2882 136715
rect 3374 65517 3434 358395
rect 3555 319292 3621 319293
rect 3555 319228 3556 319292
rect 3620 319228 3621 319292
rect 3555 319227 3621 319228
rect 3558 271829 3618 319227
rect 3739 306236 3805 306237
rect 3739 306172 3740 306236
rect 3804 306172 3805 306236
rect 3739 306171 3805 306172
rect 3555 271828 3621 271829
rect 3555 271764 3556 271828
rect 3620 271764 3621 271828
rect 3555 271763 3621 271764
rect 3555 267204 3621 267205
rect 3555 267140 3556 267204
rect 3620 267140 3621 267204
rect 3555 267139 3621 267140
rect 3558 87549 3618 267139
rect 3742 242861 3802 306171
rect 3739 242860 3805 242861
rect 3739 242796 3740 242860
rect 3804 242796 3805 242860
rect 3739 242795 3805 242796
rect 3739 162892 3805 162893
rect 3739 162828 3740 162892
rect 3804 162828 3805 162892
rect 3739 162827 3805 162828
rect 3555 87548 3621 87549
rect 3555 87484 3556 87548
rect 3620 87484 3621 87548
rect 3555 87483 3621 87484
rect 3742 76533 3802 162827
rect 3739 76532 3805 76533
rect 3739 76468 3740 76532
rect 3804 76468 3805 76532
rect 3739 76467 3805 76468
rect 4662 72453 4722 579939
rect 7419 566948 7485 566949
rect 7419 566884 7420 566948
rect 7484 566884 7485 566948
rect 7419 566883 7485 566884
rect 4843 553892 4909 553893
rect 4843 553828 4844 553892
rect 4908 553828 4909 553892
rect 4843 553827 4909 553828
rect 4846 86189 4906 553827
rect 6131 514860 6197 514861
rect 6131 514796 6132 514860
rect 6196 514796 6197 514860
rect 6131 514795 6197 514796
rect 5027 271828 5093 271829
rect 5027 271764 5028 271828
rect 5092 271764 5093 271828
rect 5027 271763 5093 271764
rect 4843 86188 4909 86189
rect 4843 86124 4844 86188
rect 4908 86124 4909 86188
rect 4843 86123 4909 86124
rect 4659 72452 4725 72453
rect 4659 72388 4660 72452
rect 4724 72388 4725 72452
rect 4659 72387 4725 72388
rect 3555 71636 3621 71637
rect 3555 71572 3556 71636
rect 3620 71572 3621 71636
rect 3555 71571 3621 71572
rect 3371 65516 3437 65517
rect 3371 65452 3372 65516
rect 3436 65452 3437 65516
rect 3371 65451 3437 65452
rect 2819 45524 2885 45525
rect 2819 45460 2820 45524
rect 2884 45460 2885 45524
rect 2819 45459 2885 45460
rect 2822 44845 2882 45459
rect 2819 44844 2885 44845
rect 2819 44780 2820 44844
rect 2884 44780 2885 44844
rect 2819 44779 2885 44780
rect 3558 22677 3618 71571
rect 3555 22676 3621 22677
rect 3555 22612 3556 22676
rect 3620 22612 3621 22676
rect 3555 22611 3621 22612
rect 2083 21724 2149 21725
rect 2083 21660 2084 21724
rect 2148 21660 2149 21724
rect 2083 21659 2149 21660
rect 243 20364 309 20365
rect 243 20300 244 20364
rect 308 20300 309 20364
rect 243 20299 309 20300
rect 5030 19005 5090 271763
rect 6134 82109 6194 514795
rect 6315 449580 6381 449581
rect 6315 449516 6316 449580
rect 6380 449516 6381 449580
rect 6315 449515 6381 449516
rect 6318 83469 6378 449515
rect 6499 397492 6565 397493
rect 6499 397428 6500 397492
rect 6564 397428 6565 397492
rect 6499 397427 6565 397428
rect 6315 83468 6381 83469
rect 6315 83404 6316 83468
rect 6380 83404 6381 83468
rect 6315 83403 6381 83404
rect 6131 82108 6197 82109
rect 6131 82044 6132 82108
rect 6196 82044 6197 82108
rect 6131 82043 6197 82044
rect 6502 77893 6562 397427
rect 7422 80749 7482 566883
rect 7603 501804 7669 501805
rect 7603 501740 7604 501804
rect 7668 501740 7669 501804
rect 7603 501739 7669 501740
rect 7606 84829 7666 501739
rect 7787 475692 7853 475693
rect 7787 475628 7788 475692
rect 7852 475628 7853 475692
rect 7787 475627 7853 475628
rect 7603 84828 7669 84829
rect 7603 84764 7604 84828
rect 7668 84764 7669 84828
rect 7603 84763 7669 84764
rect 7419 80748 7485 80749
rect 7419 80684 7420 80748
rect 7484 80684 7485 80748
rect 7419 80683 7485 80684
rect 6499 77892 6565 77893
rect 6499 77828 6500 77892
rect 6564 77828 6565 77892
rect 6499 77827 6565 77828
rect 7790 75173 7850 475627
rect 7787 75172 7853 75173
rect 7787 75108 7788 75172
rect 7852 75108 7853 75172
rect 7787 75107 7853 75108
rect 8894 69597 8954 684251
rect 285627 671260 285693 671261
rect 285627 671196 285628 671260
rect 285692 671196 285693 671260
rect 285627 671195 285693 671196
rect 281027 619172 281093 619173
rect 281027 619108 281028 619172
rect 281092 619108 281093 619172
rect 281027 619107 281093 619108
rect 9075 527916 9141 527917
rect 9075 527852 9076 527916
rect 9140 527852 9141 527916
rect 9075 527851 9141 527852
rect 9078 73813 9138 527851
rect 12387 462636 12453 462637
rect 12387 462572 12388 462636
rect 12452 462572 12453 462636
rect 12387 462571 12453 462572
rect 9259 423604 9325 423605
rect 9259 423540 9260 423604
rect 9324 423540 9325 423604
rect 9259 423539 9325 423540
rect 9262 89045 9322 423539
rect 11099 410548 11165 410549
rect 11099 410484 11100 410548
rect 11164 410484 11165 410548
rect 11099 410483 11165 410484
rect 9811 371380 9877 371381
rect 9811 371316 9812 371380
rect 9876 371316 9877 371380
rect 9811 371315 9877 371316
rect 9443 242860 9509 242861
rect 9443 242796 9444 242860
rect 9508 242796 9509 242860
rect 9443 242795 9509 242796
rect 9259 89044 9325 89045
rect 9259 88980 9260 89044
rect 9324 88980 9325 89044
rect 9259 88979 9325 88980
rect 9075 73812 9141 73813
rect 9075 73748 9076 73812
rect 9140 73748 9141 73812
rect 9075 73747 9141 73748
rect 8891 69596 8957 69597
rect 8891 69532 8892 69596
rect 8956 69532 8957 69596
rect 8891 69531 8957 69532
rect 9446 21861 9506 242795
rect 9814 200130 9874 371315
rect 10179 213892 10245 213893
rect 10179 213828 10180 213892
rect 10244 213828 10245 213892
rect 10179 213827 10245 213828
rect 9630 200070 9874 200130
rect 9630 190365 9690 200070
rect 10182 191045 10242 213827
rect 11102 213213 11162 410483
rect 12390 213893 12450 462571
rect 81672 277927 81992 278032
rect 81672 277691 81714 277927
rect 81950 277691 81992 277927
rect 81672 277586 81992 277691
rect 112392 277927 112712 278032
rect 112392 277691 112434 277927
rect 112670 277691 112712 277927
rect 112392 277586 112712 277691
rect 143112 277927 143432 278032
rect 143112 277691 143154 277927
rect 143390 277691 143432 277927
rect 143112 277586 143432 277691
rect 149936 277927 150256 278032
rect 149936 277691 149978 277927
rect 150214 277691 150256 277927
rect 149936 277586 150256 277691
rect 180656 277927 180976 278032
rect 180656 277691 180698 277927
rect 180934 277691 180976 277927
rect 180656 277586 180976 277691
rect 211376 277927 211696 278032
rect 211376 277691 211418 277927
rect 211654 277691 211696 277927
rect 211376 277586 211696 277691
rect 97032 274454 97352 274486
rect 97032 274218 97074 274454
rect 97310 274218 97352 274454
rect 97032 274134 97352 274218
rect 97032 273898 97074 274134
rect 97310 273898 97352 274134
rect 97032 273866 97352 273898
rect 127752 274454 128072 274486
rect 127752 274218 127794 274454
rect 128030 274218 128072 274454
rect 127752 274134 128072 274218
rect 127752 273898 127794 274134
rect 128030 273898 128072 274134
rect 127752 273866 128072 273898
rect 165296 274454 165616 274486
rect 165296 274218 165338 274454
rect 165574 274218 165616 274454
rect 165296 274134 165616 274218
rect 165296 273898 165338 274134
rect 165574 273898 165616 274134
rect 165296 273866 165616 273898
rect 196016 274454 196336 274486
rect 196016 274218 196058 274454
rect 196294 274218 196336 274454
rect 196016 274134 196336 274218
rect 196016 273898 196058 274134
rect 196294 273898 196336 274134
rect 196016 273866 196336 273898
rect 81672 268174 81992 268206
rect 81672 267938 81714 268174
rect 81950 267938 81992 268174
rect 81672 267854 81992 267938
rect 81672 267618 81714 267854
rect 81950 267618 81992 267854
rect 81672 267586 81992 267618
rect 112392 268174 112712 268206
rect 112392 267938 112434 268174
rect 112670 267938 112712 268174
rect 112392 267854 112712 267938
rect 112392 267618 112434 267854
rect 112670 267618 112712 267854
rect 112392 267586 112712 267618
rect 143112 268174 143432 268206
rect 143112 267938 143154 268174
rect 143390 267938 143432 268174
rect 143112 267854 143432 267938
rect 143112 267618 143154 267854
rect 143390 267618 143432 267854
rect 143112 267586 143432 267618
rect 149936 268174 150256 268206
rect 149936 267938 149978 268174
rect 150214 267938 150256 268174
rect 149936 267854 150256 267938
rect 149936 267618 149978 267854
rect 150214 267618 150256 267854
rect 149936 267586 150256 267618
rect 180656 268174 180976 268206
rect 180656 267938 180698 268174
rect 180934 267938 180976 268174
rect 180656 267854 180976 267938
rect 180656 267618 180698 267854
rect 180934 267618 180976 267854
rect 180656 267586 180976 267618
rect 211376 268174 211696 268206
rect 211376 267938 211418 268174
rect 211654 267938 211696 268174
rect 211376 267854 211696 267938
rect 211376 267618 211418 267854
rect 211654 267618 211696 267854
rect 211376 267586 211696 267618
rect 97032 264454 97352 264486
rect 97032 264218 97074 264454
rect 97310 264218 97352 264454
rect 97032 264134 97352 264218
rect 97032 263898 97074 264134
rect 97310 263898 97352 264134
rect 97032 263866 97352 263898
rect 127752 264454 128072 264486
rect 127752 264218 127794 264454
rect 128030 264218 128072 264454
rect 127752 264134 128072 264218
rect 127752 263898 127794 264134
rect 128030 263898 128072 264134
rect 127752 263866 128072 263898
rect 165296 264454 165616 264486
rect 165296 264218 165338 264454
rect 165574 264218 165616 264454
rect 165296 264134 165616 264218
rect 165296 263898 165338 264134
rect 165574 263898 165616 264134
rect 165296 263866 165616 263898
rect 196016 264454 196336 264486
rect 196016 264218 196058 264454
rect 196294 264218 196336 264454
rect 196016 264134 196336 264218
rect 196016 263898 196058 264134
rect 196294 263898 196336 264134
rect 196016 263866 196336 263898
rect 81672 258174 81992 258206
rect 81672 257938 81714 258174
rect 81950 257938 81992 258174
rect 81672 257854 81992 257938
rect 81672 257618 81714 257854
rect 81950 257618 81992 257854
rect 81672 257586 81992 257618
rect 112392 258174 112712 258206
rect 112392 257938 112434 258174
rect 112670 257938 112712 258174
rect 112392 257854 112712 257938
rect 112392 257618 112434 257854
rect 112670 257618 112712 257854
rect 112392 257586 112712 257618
rect 143112 258174 143432 258206
rect 143112 257938 143154 258174
rect 143390 257938 143432 258174
rect 143112 257854 143432 257938
rect 143112 257618 143154 257854
rect 143390 257618 143432 257854
rect 143112 257586 143432 257618
rect 149936 258174 150256 258206
rect 149936 257938 149978 258174
rect 150214 257938 150256 258174
rect 149936 257854 150256 257938
rect 149936 257618 149978 257854
rect 150214 257618 150256 257854
rect 149936 257586 150256 257618
rect 180656 258174 180976 258206
rect 180656 257938 180698 258174
rect 180934 257938 180976 258174
rect 180656 257854 180976 257938
rect 180656 257618 180698 257854
rect 180934 257618 180976 257854
rect 180656 257586 180976 257618
rect 211376 258174 211696 258206
rect 211376 257938 211418 258174
rect 211654 257938 211696 258174
rect 211376 257854 211696 257938
rect 211376 257618 211418 257854
rect 211654 257618 211696 257854
rect 211376 257586 211696 257618
rect 97032 254454 97352 254486
rect 97032 254218 97074 254454
rect 97310 254218 97352 254454
rect 97032 254134 97352 254218
rect 97032 253898 97074 254134
rect 97310 253898 97352 254134
rect 97032 253866 97352 253898
rect 127752 254454 128072 254486
rect 127752 254218 127794 254454
rect 128030 254218 128072 254454
rect 127752 254134 128072 254218
rect 127752 253898 127794 254134
rect 128030 253898 128072 254134
rect 127752 253866 128072 253898
rect 165296 254454 165616 254486
rect 165296 254218 165338 254454
rect 165574 254218 165616 254454
rect 165296 254134 165616 254218
rect 165296 253898 165338 254134
rect 165574 253898 165616 254134
rect 165296 253866 165616 253898
rect 196016 254454 196336 254486
rect 196016 254218 196058 254454
rect 196294 254218 196336 254454
rect 196016 254134 196336 254218
rect 196016 253898 196058 254134
rect 196294 253898 196336 254134
rect 196016 253866 196336 253898
rect 81672 248174 81992 248206
rect 81672 247938 81714 248174
rect 81950 247938 81992 248174
rect 81672 247854 81992 247938
rect 81672 247618 81714 247854
rect 81950 247618 81992 247854
rect 81672 247586 81992 247618
rect 112392 248174 112712 248206
rect 112392 247938 112434 248174
rect 112670 247938 112712 248174
rect 112392 247854 112712 247938
rect 112392 247618 112434 247854
rect 112670 247618 112712 247854
rect 112392 247586 112712 247618
rect 143112 248174 143432 248206
rect 143112 247938 143154 248174
rect 143390 247938 143432 248174
rect 143112 247854 143432 247938
rect 143112 247618 143154 247854
rect 143390 247618 143432 247854
rect 143112 247586 143432 247618
rect 149936 248174 150256 248206
rect 149936 247938 149978 248174
rect 150214 247938 150256 248174
rect 149936 247854 150256 247938
rect 149936 247618 149978 247854
rect 150214 247618 150256 247854
rect 149936 247586 150256 247618
rect 180656 248174 180976 248206
rect 180656 247938 180698 248174
rect 180934 247938 180976 248174
rect 180656 247854 180976 247938
rect 180656 247618 180698 247854
rect 180934 247618 180976 247854
rect 180656 247586 180976 247618
rect 211376 248174 211696 248206
rect 211376 247938 211418 248174
rect 211654 247938 211696 248174
rect 211376 247854 211696 247938
rect 211376 247618 211418 247854
rect 211654 247618 211696 247854
rect 211376 247586 211696 247618
rect 97032 244454 97352 244486
rect 97032 244218 97074 244454
rect 97310 244218 97352 244454
rect 97032 244134 97352 244218
rect 97032 243898 97074 244134
rect 97310 243898 97352 244134
rect 97032 243866 97352 243898
rect 127752 244454 128072 244486
rect 127752 244218 127794 244454
rect 128030 244218 128072 244454
rect 127752 244134 128072 244218
rect 127752 243898 127794 244134
rect 128030 243898 128072 244134
rect 127752 243866 128072 243898
rect 165296 244454 165616 244486
rect 165296 244218 165338 244454
rect 165574 244218 165616 244454
rect 165296 244134 165616 244218
rect 165296 243898 165338 244134
rect 165574 243898 165616 244134
rect 165296 243866 165616 243898
rect 196016 244454 196336 244486
rect 196016 244218 196058 244454
rect 196294 244218 196336 244454
rect 196016 244134 196336 244218
rect 196016 243898 196058 244134
rect 196294 243898 196336 244134
rect 196016 243866 196336 243898
rect 81672 238174 81992 238206
rect 81672 237938 81714 238174
rect 81950 237938 81992 238174
rect 81672 237854 81992 237938
rect 81672 237618 81714 237854
rect 81950 237618 81992 237854
rect 81672 237586 81992 237618
rect 112392 238174 112712 238206
rect 112392 237938 112434 238174
rect 112670 237938 112712 238174
rect 112392 237854 112712 237938
rect 112392 237618 112434 237854
rect 112670 237618 112712 237854
rect 112392 237586 112712 237618
rect 143112 238174 143432 238206
rect 143112 237938 143154 238174
rect 143390 237938 143432 238174
rect 143112 237854 143432 237938
rect 143112 237618 143154 237854
rect 143390 237618 143432 237854
rect 143112 237586 143432 237618
rect 149936 238174 150256 238206
rect 149936 237938 149978 238174
rect 150214 237938 150256 238174
rect 149936 237854 150256 237938
rect 149936 237618 149978 237854
rect 150214 237618 150256 237854
rect 149936 237586 150256 237618
rect 180656 238174 180976 238206
rect 180656 237938 180698 238174
rect 180934 237938 180976 238174
rect 180656 237854 180976 237938
rect 180656 237618 180698 237854
rect 180934 237618 180976 237854
rect 180656 237586 180976 237618
rect 211376 238174 211696 238206
rect 211376 237938 211418 238174
rect 211654 237938 211696 238174
rect 211376 237854 211696 237938
rect 211376 237618 211418 237854
rect 211654 237618 211696 237854
rect 211376 237586 211696 237618
rect 78443 234020 78509 234021
rect 78443 233956 78444 234020
rect 78508 233956 78509 234020
rect 78443 233955 78509 233956
rect 12387 213892 12453 213893
rect 12387 213828 12388 213892
rect 12452 213828 12453 213892
rect 12387 213827 12453 213828
rect 11099 213212 11165 213213
rect 11099 213148 11100 213212
rect 11164 213148 11165 213212
rect 11099 213147 11165 213148
rect 14065 208174 14385 208206
rect 14065 207938 14107 208174
rect 14343 207938 14385 208174
rect 14065 207854 14385 207938
rect 14065 207618 14107 207854
rect 14343 207618 14385 207854
rect 14065 207586 14385 207618
rect 21907 208174 22227 208206
rect 21907 207938 21949 208174
rect 22185 207938 22227 208174
rect 21907 207854 22227 207938
rect 21907 207618 21949 207854
rect 22185 207618 22227 207854
rect 21907 207586 22227 207618
rect 29749 208174 30069 208206
rect 29749 207938 29791 208174
rect 30027 207938 30069 208174
rect 29749 207854 30069 207938
rect 29749 207618 29791 207854
rect 30027 207618 30069 207854
rect 29749 207586 30069 207618
rect 37591 208174 37911 208206
rect 37591 207938 37633 208174
rect 37869 207938 37911 208174
rect 37591 207854 37911 207938
rect 37591 207618 37633 207854
rect 37869 207618 37911 207854
rect 37591 207586 37911 207618
rect 42248 208174 43248 208206
rect 42248 207938 42310 208174
rect 42546 207938 42630 208174
rect 42866 207938 42950 208174
rect 43186 207938 43248 208174
rect 42248 207854 43248 207938
rect 42248 207618 42310 207854
rect 42546 207618 42630 207854
rect 42866 207618 42950 207854
rect 43186 207618 43248 207854
rect 42248 207586 43248 207618
rect 17986 204454 18306 204486
rect 17986 204218 18028 204454
rect 18264 204218 18306 204454
rect 17986 204134 18306 204218
rect 17986 203898 18028 204134
rect 18264 203898 18306 204134
rect 17986 203866 18306 203898
rect 25828 204454 26148 204486
rect 25828 204218 25870 204454
rect 26106 204218 26148 204454
rect 25828 204134 26148 204218
rect 25828 203898 25870 204134
rect 26106 203898 26148 204134
rect 25828 203866 26148 203898
rect 33670 204454 33990 204486
rect 33670 204218 33712 204454
rect 33948 204218 33990 204454
rect 33670 204134 33990 204218
rect 33670 203898 33712 204134
rect 33948 203898 33990 204134
rect 33670 203866 33990 203898
rect 41512 204454 41832 204486
rect 41512 204218 41554 204454
rect 41790 204218 41832 204454
rect 41512 204134 41832 204218
rect 41512 203898 41554 204134
rect 41790 203898 41832 204134
rect 41512 203866 41832 203898
rect 52118 204454 52438 204486
rect 52118 204218 52160 204454
rect 52396 204218 52438 204454
rect 52118 204134 52438 204218
rect 52118 203898 52160 204134
rect 52396 203898 52438 204134
rect 52118 203866 52438 203898
rect 59960 204454 60280 204486
rect 59960 204218 60002 204454
rect 60238 204218 60280 204454
rect 59960 204134 60280 204218
rect 59960 203898 60002 204134
rect 60238 203898 60280 204134
rect 59960 203866 60280 203898
rect 67802 204454 68122 204486
rect 67802 204218 67844 204454
rect 68080 204218 68122 204454
rect 67802 204134 68122 204218
rect 67802 203898 67844 204134
rect 68080 203898 68122 204134
rect 67802 203866 68122 203898
rect 75644 204454 75964 204486
rect 75644 204218 75686 204454
rect 75922 204218 75964 204454
rect 75644 204134 75964 204218
rect 75644 203898 75686 204134
rect 75922 203898 75964 204134
rect 75644 203866 75964 203898
rect 14065 198174 14385 198206
rect 14065 197938 14107 198174
rect 14343 197938 14385 198174
rect 14065 197854 14385 197938
rect 14065 197618 14107 197854
rect 14343 197618 14385 197854
rect 14065 197586 14385 197618
rect 21907 198174 22227 198206
rect 21907 197938 21949 198174
rect 22185 197938 22227 198174
rect 21907 197854 22227 197938
rect 21907 197618 21949 197854
rect 22185 197618 22227 197854
rect 21907 197586 22227 197618
rect 29749 198174 30069 198206
rect 29749 197938 29791 198174
rect 30027 197938 30069 198174
rect 29749 197854 30069 197938
rect 29749 197618 29791 197854
rect 30027 197618 30069 197854
rect 29749 197586 30069 197618
rect 37591 198174 37911 198206
rect 37591 197938 37633 198174
rect 37869 197938 37911 198174
rect 37591 197854 37911 197938
rect 37591 197618 37633 197854
rect 37869 197618 37911 197854
rect 37591 197586 37911 197618
rect 42248 198174 43248 198206
rect 42248 197938 42310 198174
rect 42546 197938 42630 198174
rect 42866 197938 42950 198174
rect 43186 197938 43248 198174
rect 42248 197854 43248 197938
rect 42248 197618 42310 197854
rect 42546 197618 42630 197854
rect 42866 197618 42950 197854
rect 43186 197618 43248 197854
rect 42248 197586 43248 197618
rect 17986 194454 18306 194486
rect 17986 194218 18028 194454
rect 18264 194218 18306 194454
rect 17986 194134 18306 194218
rect 17986 193898 18028 194134
rect 18264 193898 18306 194134
rect 17986 193866 18306 193898
rect 25828 194454 26148 194486
rect 25828 194218 25870 194454
rect 26106 194218 26148 194454
rect 25828 194134 26148 194218
rect 25828 193898 25870 194134
rect 26106 193898 26148 194134
rect 25828 193866 26148 193898
rect 33670 194454 33990 194486
rect 33670 194218 33712 194454
rect 33948 194218 33990 194454
rect 33670 194134 33990 194218
rect 33670 193898 33712 194134
rect 33948 193898 33990 194134
rect 33670 193866 33990 193898
rect 41512 194454 41832 194486
rect 41512 194218 41554 194454
rect 41790 194218 41832 194454
rect 41512 194134 41832 194218
rect 41512 193898 41554 194134
rect 41790 193898 41832 194134
rect 41512 193866 41832 193898
rect 52118 194454 52438 194486
rect 52118 194218 52160 194454
rect 52396 194218 52438 194454
rect 52118 194134 52438 194218
rect 52118 193898 52160 194134
rect 52396 193898 52438 194134
rect 52118 193866 52438 193898
rect 59960 194454 60280 194486
rect 59960 194218 60002 194454
rect 60238 194218 60280 194454
rect 59960 194134 60280 194218
rect 59960 193898 60002 194134
rect 60238 193898 60280 194134
rect 59960 193866 60280 193898
rect 67802 194454 68122 194486
rect 67802 194218 67844 194454
rect 68080 194218 68122 194454
rect 67802 194134 68122 194218
rect 67802 193898 67844 194134
rect 68080 193898 68122 194134
rect 67802 193866 68122 193898
rect 75644 194454 75964 194486
rect 75644 194218 75686 194454
rect 75922 194218 75964 194454
rect 75644 194134 75964 194218
rect 75644 193898 75686 194134
rect 75922 193898 75964 194134
rect 75644 193866 75964 193898
rect 78446 192677 78506 233955
rect 78443 192676 78509 192677
rect 78443 192612 78444 192676
rect 78508 192612 78509 192676
rect 78443 192611 78509 192612
rect 10179 191044 10245 191045
rect 10179 190980 10180 191044
rect 10244 190980 10245 191044
rect 10179 190979 10245 190980
rect 10734 190400 10794 191080
rect 11470 190400 11530 191080
rect 12206 190400 12266 191080
rect 12942 190400 13002 191080
rect 13678 190400 13738 191080
rect 14414 190400 14474 191080
rect 15150 190400 15210 191080
rect 15886 190400 15946 191080
rect 16622 190400 16682 191080
rect 17358 190400 17418 191080
rect 18094 190400 18154 191080
rect 18830 190400 18890 191080
rect 19566 190400 19626 191080
rect 20302 190400 20362 191080
rect 21038 190400 21098 191080
rect 21774 190400 21834 191080
rect 22510 190400 22570 191080
rect 23246 190400 23306 191080
rect 23982 190400 24042 191080
rect 24718 190400 24778 191080
rect 25454 190400 25514 191080
rect 26190 190400 26250 191080
rect 26926 190400 26986 191080
rect 27662 190400 27722 191080
rect 9627 190364 9693 190365
rect 9627 190300 9628 190364
rect 9692 190300 9693 190364
rect 9627 190299 9693 190300
rect 28398 190060 28458 191044
rect 29134 190400 29194 191044
rect 29870 190060 29930 191044
rect 30606 190060 30666 191044
rect 31342 190060 31402 191044
rect 32078 190060 32138 191044
rect 32814 190060 32874 191044
rect 33550 190400 33610 191044
rect 34286 190060 34346 191080
rect 35022 190400 35082 191080
rect 35758 190400 35818 191080
rect 36494 190060 36554 191080
rect 37230 190060 37290 191044
rect 37966 190060 38026 191044
rect 38702 190400 38762 191044
rect 39438 190400 39498 191080
rect 40174 190060 40234 191044
rect 40910 190400 40970 191044
rect 41646 190400 41706 191044
rect 44866 190770 44926 191420
rect 44774 190710 44926 190770
rect 44774 190470 44834 190710
rect 44774 190410 44926 190470
rect 44866 190400 44926 190410
rect 45602 190400 45662 191080
rect 46338 190400 46398 191080
rect 47074 190770 47134 191420
rect 46982 190710 47134 190770
rect 46982 190470 47042 190710
rect 46982 190410 47134 190470
rect 47074 190400 47134 190410
rect 47810 190400 47870 191080
rect 48546 190400 48606 191080
rect 49282 190400 49342 191080
rect 50018 190400 50078 191080
rect 50754 190400 50814 191080
rect 51490 190400 51550 191080
rect 52226 190400 52286 191080
rect 52962 190400 53022 191420
rect 53698 190400 53758 191080
rect 54434 190400 54494 191080
rect 55170 190400 55230 191080
rect 55906 190400 55966 191080
rect 56642 190400 56702 191080
rect 57378 190400 57438 191080
rect 58114 190400 58174 191080
rect 58850 190400 58910 191080
rect 59586 190400 59646 191080
rect 60322 190400 60382 191080
rect 61058 190400 61118 191080
rect 61794 190400 61854 191080
rect 62530 190400 62590 191080
rect 63266 190400 63326 191080
rect 64002 190400 64062 191080
rect 64738 190400 64798 191080
rect 65474 190400 65534 191080
rect 66210 190400 66270 191080
rect 66946 190400 67006 191080
rect 67682 190400 67742 191080
rect 68418 190400 68478 191044
rect 69154 190400 69214 191044
rect 69890 190400 69950 191044
rect 70626 190400 70686 191044
rect 71362 190400 71422 191044
rect 72098 190400 72158 191044
rect 72834 190400 72894 191044
rect 73570 190400 73630 191080
rect 74306 190400 74366 191080
rect 75042 190400 75102 191080
rect 75778 190400 75838 191044
rect 78998 190400 79058 235620
rect 79734 190400 79794 235162
rect 80470 190400 80530 235620
rect 81206 190400 81266 235620
rect 81942 190400 82002 235280
rect 82678 190060 82738 235620
rect 83414 190400 83474 235620
rect 84150 234970 84210 235620
rect 83966 234910 84210 234970
rect 83966 190470 84026 234910
rect 83966 190410 84210 190470
rect 84150 190060 84210 190410
rect 84886 190400 84946 235162
rect 85622 190400 85682 235162
rect 86358 190400 86418 235162
rect 87094 190400 87154 235280
rect 87830 190400 87890 235620
rect 88566 190400 88626 235620
rect 89302 233885 89362 235620
rect 90038 234021 90098 235620
rect 90035 234020 90101 234021
rect 90035 233956 90036 234020
rect 90100 233956 90101 234020
rect 90035 233955 90101 233956
rect 89299 233884 89365 233885
rect 89299 233820 89300 233884
rect 89364 233820 89365 233884
rect 89299 233819 89365 233820
rect 90035 192676 90101 192677
rect 90035 192612 90036 192676
rect 90100 192612 90101 192676
rect 90035 192611 90101 192612
rect 89299 192540 89365 192541
rect 89299 192476 89300 192540
rect 89364 192476 89365 192540
rect 89299 192475 89365 192476
rect 89302 190400 89362 192475
rect 90038 190400 90098 192611
rect 90774 190400 90834 235620
rect 91510 190400 91570 235280
rect 92246 190400 92306 235162
rect 92982 190400 93042 235620
rect 93718 190400 93778 235162
rect 94454 190400 94514 235162
rect 95190 190400 95250 235162
rect 95926 190400 95986 235162
rect 96662 190060 96722 235108
rect 97398 190400 97458 235108
rect 98134 190060 98194 235108
rect 98870 190400 98930 235108
rect 99606 190060 99666 235108
rect 100342 190400 100402 235108
rect 101078 190400 101138 235108
rect 101814 190400 101874 235108
rect 102550 190400 102610 235108
rect 103286 190060 103346 235108
rect 104022 190060 104082 235620
rect 104758 190400 104818 235162
rect 105494 190400 105554 235280
rect 106230 229110 106290 235162
rect 106230 229050 106474 229110
rect 106414 190470 106474 229050
rect 106230 190410 106474 190470
rect 106230 190060 106290 190410
rect 106966 190060 107026 235280
rect 107702 190400 107762 235162
rect 108438 190060 108498 235162
rect 109174 190400 109234 235125
rect 109910 190400 109970 235108
rect 110459 233884 110525 233885
rect 110459 233820 110460 233884
rect 110524 233820 110525 233884
rect 110459 233819 110525 233820
rect 110462 192541 110522 233819
rect 116461 228174 116781 228206
rect 116461 227938 116503 228174
rect 116739 227938 116781 228174
rect 116461 227854 116781 227938
rect 116461 227618 116503 227854
rect 116739 227618 116781 227854
rect 116461 227586 116781 227618
rect 124303 228174 124623 228206
rect 124303 227938 124345 228174
rect 124581 227938 124623 228174
rect 124303 227854 124623 227938
rect 124303 227618 124345 227854
rect 124581 227618 124623 227854
rect 124303 227586 124623 227618
rect 132145 228174 132465 228206
rect 132145 227938 132187 228174
rect 132423 227938 132465 228174
rect 132145 227854 132465 227938
rect 132145 227618 132187 227854
rect 132423 227618 132465 227854
rect 132145 227586 132465 227618
rect 139987 228174 140307 228206
rect 139987 227938 140029 228174
rect 140265 227938 140307 228174
rect 139987 227854 140307 227938
rect 139987 227618 140029 227854
rect 140265 227618 140307 227854
rect 139987 227586 140307 227618
rect 120382 224454 120702 224486
rect 120382 224218 120424 224454
rect 120660 224218 120702 224454
rect 120382 224134 120702 224218
rect 120382 223898 120424 224134
rect 120660 223898 120702 224134
rect 120382 223866 120702 223898
rect 128224 224454 128544 224486
rect 128224 224218 128266 224454
rect 128502 224218 128544 224454
rect 128224 224134 128544 224218
rect 128224 223898 128266 224134
rect 128502 223898 128544 224134
rect 128224 223866 128544 223898
rect 136066 224454 136386 224486
rect 136066 224218 136108 224454
rect 136344 224218 136386 224454
rect 136066 224134 136386 224218
rect 136066 223898 136108 224134
rect 136344 223898 136386 224134
rect 136066 223866 136386 223898
rect 143908 224454 144228 224486
rect 143908 224218 143950 224454
rect 144186 224218 144228 224454
rect 143908 224134 144228 224218
rect 143908 223898 143950 224134
rect 144186 223898 144228 224134
rect 143908 223866 144228 223898
rect 116461 218174 116781 218206
rect 116461 217938 116503 218174
rect 116739 217938 116781 218174
rect 116461 217854 116781 217938
rect 116461 217618 116503 217854
rect 116739 217618 116781 217854
rect 116461 217586 116781 217618
rect 124303 218174 124623 218206
rect 124303 217938 124345 218174
rect 124581 217938 124623 218174
rect 124303 217854 124623 217938
rect 124303 217618 124345 217854
rect 124581 217618 124623 217854
rect 124303 217586 124623 217618
rect 132145 218174 132465 218206
rect 132145 217938 132187 218174
rect 132423 217938 132465 218174
rect 132145 217854 132465 217938
rect 132145 217618 132187 217854
rect 132423 217618 132465 217854
rect 132145 217586 132465 217618
rect 139987 218174 140307 218206
rect 139987 217938 140029 218174
rect 140265 217938 140307 218174
rect 139987 217854 140307 217938
rect 139987 217618 140029 217854
rect 140265 217618 140307 217854
rect 139987 217586 140307 217618
rect 120382 214454 120702 214486
rect 120382 214218 120424 214454
rect 120660 214218 120702 214454
rect 120382 214134 120702 214218
rect 120382 213898 120424 214134
rect 120660 213898 120702 214134
rect 120382 213866 120702 213898
rect 128224 214454 128544 214486
rect 128224 214218 128266 214454
rect 128502 214218 128544 214454
rect 128224 214134 128544 214218
rect 128224 213898 128266 214134
rect 128502 213898 128544 214134
rect 128224 213866 128544 213898
rect 136066 214454 136386 214486
rect 136066 214218 136108 214454
rect 136344 214218 136386 214454
rect 136066 214134 136386 214218
rect 136066 213898 136108 214134
rect 136344 213898 136386 214134
rect 136066 213866 136386 213898
rect 143908 214454 144228 214486
rect 143908 214218 143950 214454
rect 144186 214218 144228 214454
rect 143908 214134 144228 214218
rect 143908 213898 143950 214134
rect 144186 213898 144228 214134
rect 143908 213866 144228 213898
rect 116461 208174 116781 208206
rect 116461 207938 116503 208174
rect 116739 207938 116781 208174
rect 116461 207854 116781 207938
rect 116461 207618 116503 207854
rect 116739 207618 116781 207854
rect 116461 207586 116781 207618
rect 124303 208174 124623 208206
rect 124303 207938 124345 208174
rect 124581 207938 124623 208174
rect 124303 207854 124623 207938
rect 124303 207618 124345 207854
rect 124581 207618 124623 207854
rect 124303 207586 124623 207618
rect 132145 208174 132465 208206
rect 132145 207938 132187 208174
rect 132423 207938 132465 208174
rect 132145 207854 132465 207938
rect 132145 207618 132187 207854
rect 132423 207618 132465 207854
rect 132145 207586 132465 207618
rect 139987 208174 140307 208206
rect 139987 207938 140029 208174
rect 140265 207938 140307 208174
rect 139987 207854 140307 207938
rect 139987 207618 140029 207854
rect 140265 207618 140307 207854
rect 139987 207586 140307 207618
rect 120382 204454 120702 204486
rect 120382 204218 120424 204454
rect 120660 204218 120702 204454
rect 120382 204134 120702 204218
rect 120382 203898 120424 204134
rect 120660 203898 120702 204134
rect 120382 203866 120702 203898
rect 128224 204454 128544 204486
rect 128224 204218 128266 204454
rect 128502 204218 128544 204454
rect 128224 204134 128544 204218
rect 128224 203898 128266 204134
rect 128502 203898 128544 204134
rect 128224 203866 128544 203898
rect 136066 204454 136386 204486
rect 136066 204218 136108 204454
rect 136344 204218 136386 204454
rect 136066 204134 136386 204218
rect 136066 203898 136108 204134
rect 136344 203898 136386 204134
rect 136066 203866 136386 203898
rect 143908 204454 144228 204486
rect 143908 204218 143950 204454
rect 144186 204218 144228 204454
rect 143908 204134 144228 204218
rect 143908 203898 143950 204134
rect 144186 203898 144228 204134
rect 143908 203866 144228 203898
rect 116461 198174 116781 198206
rect 116461 197938 116503 198174
rect 116739 197938 116781 198174
rect 116461 197854 116781 197938
rect 116461 197618 116503 197854
rect 116739 197618 116781 197854
rect 116461 197586 116781 197618
rect 124303 198174 124623 198206
rect 124303 197938 124345 198174
rect 124581 197938 124623 198174
rect 124303 197854 124623 197938
rect 124303 197618 124345 197854
rect 124581 197618 124623 197854
rect 124303 197586 124623 197618
rect 132145 198174 132465 198206
rect 132145 197938 132187 198174
rect 132423 197938 132465 198174
rect 132145 197854 132465 197938
rect 132145 197618 132187 197854
rect 132423 197618 132465 197854
rect 132145 197586 132465 197618
rect 139987 198174 140307 198206
rect 139987 197938 140029 198174
rect 140265 197938 140307 198174
rect 139987 197854 140307 197938
rect 139987 197618 140029 197854
rect 140265 197618 140307 197854
rect 139987 197586 140307 197618
rect 120382 194454 120702 194486
rect 120382 194218 120424 194454
rect 120660 194218 120702 194454
rect 120382 194134 120702 194218
rect 120382 193898 120424 194134
rect 120660 193898 120702 194134
rect 120382 193866 120702 193898
rect 128224 194454 128544 194486
rect 128224 194218 128266 194454
rect 128502 194218 128544 194454
rect 128224 194134 128544 194218
rect 128224 193898 128266 194134
rect 128502 193898 128544 194134
rect 128224 193866 128544 193898
rect 136066 194454 136386 194486
rect 136066 194218 136108 194454
rect 136344 194218 136386 194454
rect 136066 194134 136386 194218
rect 136066 193898 136108 194134
rect 136344 193898 136386 194134
rect 136066 193866 136386 193898
rect 143908 194454 144228 194486
rect 143908 194218 143950 194454
rect 144186 194218 144228 194454
rect 143908 194134 144228 194218
rect 143908 193898 143950 194134
rect 144186 193898 144228 194134
rect 143908 193866 144228 193898
rect 110459 192540 110525 192541
rect 110459 192476 110460 192540
rect 110524 192476 110525 192540
rect 110459 192475 110525 192476
rect 113130 190400 113190 191080
rect 113866 190400 113926 191080
rect 114602 190400 114662 191080
rect 115338 190400 115398 191080
rect 116074 190400 116134 191080
rect 116810 190400 116870 191080
rect 117546 190400 117606 191080
rect 118282 190400 118342 191080
rect 119018 190400 119078 191080
rect 119754 190400 119814 191080
rect 120490 190400 120550 191080
rect 121226 190400 121286 191080
rect 121962 190400 122022 191080
rect 122698 190400 122758 191080
rect 123434 190400 123494 191080
rect 124170 190400 124230 191080
rect 124906 190400 124966 191420
rect 125642 190400 125702 191420
rect 126378 190400 126438 191420
rect 127114 190400 127174 191080
rect 127850 190400 127910 191080
rect 128586 190400 128646 191080
rect 129322 190400 129382 191420
rect 130058 190400 130118 191080
rect 130794 190400 130854 191044
rect 131530 190400 131590 191044
rect 132266 190400 132326 191044
rect 133002 190400 133062 191044
rect 133738 190400 133798 191044
rect 134474 190400 134534 191044
rect 135210 190400 135270 191044
rect 135946 190400 136006 191044
rect 136682 190400 136742 191080
rect 137418 190400 137478 191080
rect 138154 190400 138214 191080
rect 138890 190400 138950 191080
rect 139626 190400 139686 191080
rect 140362 190400 140422 191080
rect 141098 190400 141158 191080
rect 141834 190400 141894 191044
rect 142570 190400 142630 191044
rect 143306 190400 143366 191080
rect 144042 190400 144102 191044
rect 147262 190400 147322 235280
rect 147998 190400 148058 235280
rect 148734 190400 148794 235280
rect 149470 190400 149530 235280
rect 150206 190400 150266 235280
rect 150942 190400 151002 235280
rect 151678 190400 151738 235280
rect 152414 190400 152474 235280
rect 153150 190400 153210 235280
rect 153886 190400 153946 235280
rect 154622 190400 154682 235162
rect 155358 190400 155418 235162
rect 156094 190400 156154 235280
rect 156830 190400 156890 235280
rect 157566 190400 157626 235280
rect 158302 190400 158362 235162
rect 159038 190400 159098 235162
rect 159774 190400 159834 235162
rect 160510 190400 160570 235162
rect 161246 190400 161306 235280
rect 161982 190400 162042 235162
rect 162718 190400 162778 235162
rect 163454 190400 163514 235280
rect 164190 229110 164250 235280
rect 164190 229050 164434 229110
rect 164374 190470 164434 229050
rect 164190 190410 164434 190470
rect 164190 190400 164250 190410
rect 164926 190060 164986 235108
rect 165662 190400 165722 235108
rect 166398 190060 166458 235108
rect 167134 190060 167194 235108
rect 167870 190060 167930 235108
rect 168606 190060 168666 235108
rect 169342 190060 169402 235108
rect 170078 190060 170138 235108
rect 170814 190060 170874 235108
rect 171550 190060 171610 235108
rect 172286 190060 172346 235108
rect 173022 190060 173082 235108
rect 173758 190060 173818 235108
rect 174494 190060 174554 235162
rect 175230 190060 175290 235162
rect 175966 190060 176026 235230
rect 176702 190400 176762 235162
rect 177438 190400 177498 235620
rect 178174 190400 178234 235108
rect 184725 208174 185045 208206
rect 184725 207938 184767 208174
rect 185003 207938 185045 208174
rect 184725 207854 185045 207938
rect 184725 207618 184767 207854
rect 185003 207618 185045 207854
rect 184725 207586 185045 207618
rect 192567 208174 192887 208206
rect 192567 207938 192609 208174
rect 192845 207938 192887 208174
rect 192567 207854 192887 207938
rect 192567 207618 192609 207854
rect 192845 207618 192887 207854
rect 192567 207586 192887 207618
rect 200409 208174 200729 208206
rect 200409 207938 200451 208174
rect 200687 207938 200729 208174
rect 200409 207854 200729 207938
rect 200409 207618 200451 207854
rect 200687 207618 200729 207854
rect 200409 207586 200729 207618
rect 208251 208174 208571 208206
rect 208251 207938 208293 208174
rect 208529 207938 208571 208174
rect 208251 207854 208571 207938
rect 208251 207618 208293 207854
rect 208529 207618 208571 207854
rect 208251 207586 208571 207618
rect 218857 208174 219177 208206
rect 218857 207938 218899 208174
rect 219135 207938 219177 208174
rect 218857 207854 219177 207938
rect 218857 207618 218899 207854
rect 219135 207618 219177 207854
rect 218857 207586 219177 207618
rect 226699 208174 227019 208206
rect 226699 207938 226741 208174
rect 226977 207938 227019 208174
rect 226699 207854 227019 207938
rect 226699 207618 226741 207854
rect 226977 207618 227019 207854
rect 226699 207586 227019 207618
rect 234541 208174 234861 208206
rect 234541 207938 234583 208174
rect 234819 207938 234861 208174
rect 234541 207854 234861 207938
rect 234541 207618 234583 207854
rect 234819 207618 234861 207854
rect 234541 207586 234861 207618
rect 242383 208174 242703 208206
rect 242383 207938 242425 208174
rect 242661 207938 242703 208174
rect 242383 207854 242703 207938
rect 242383 207618 242425 207854
rect 242661 207618 242703 207854
rect 242383 207586 242703 207618
rect 252989 208174 253309 208206
rect 252989 207938 253031 208174
rect 253267 207938 253309 208174
rect 252989 207854 253309 207938
rect 252989 207618 253031 207854
rect 253267 207618 253309 207854
rect 252989 207586 253309 207618
rect 260831 208174 261151 208206
rect 260831 207938 260873 208174
rect 261109 207938 261151 208174
rect 260831 207854 261151 207938
rect 260831 207618 260873 207854
rect 261109 207618 261151 207854
rect 260831 207586 261151 207618
rect 268673 208174 268993 208206
rect 268673 207938 268715 208174
rect 268951 207938 268993 208174
rect 268673 207854 268993 207938
rect 268673 207618 268715 207854
rect 268951 207618 268993 207854
rect 268673 207586 268993 207618
rect 276515 208174 276835 208206
rect 276515 207938 276557 208174
rect 276793 207938 276835 208174
rect 276515 207854 276835 207938
rect 276515 207618 276557 207854
rect 276793 207618 276835 207854
rect 276515 207586 276835 207618
rect 188646 204454 188966 204486
rect 188646 204218 188688 204454
rect 188924 204218 188966 204454
rect 188646 204134 188966 204218
rect 188646 203898 188688 204134
rect 188924 203898 188966 204134
rect 188646 203866 188966 203898
rect 196488 204454 196808 204486
rect 196488 204218 196530 204454
rect 196766 204218 196808 204454
rect 196488 204134 196808 204218
rect 196488 203898 196530 204134
rect 196766 203898 196808 204134
rect 196488 203866 196808 203898
rect 204330 204454 204650 204486
rect 204330 204218 204372 204454
rect 204608 204218 204650 204454
rect 204330 204134 204650 204218
rect 204330 203898 204372 204134
rect 204608 203898 204650 204134
rect 204330 203866 204650 203898
rect 212172 204454 212492 204486
rect 212172 204218 212214 204454
rect 212450 204218 212492 204454
rect 212172 204134 212492 204218
rect 212172 203898 212214 204134
rect 212450 203898 212492 204134
rect 212172 203866 212492 203898
rect 222778 204454 223098 204486
rect 222778 204218 222820 204454
rect 223056 204218 223098 204454
rect 222778 204134 223098 204218
rect 222778 203898 222820 204134
rect 223056 203898 223098 204134
rect 222778 203866 223098 203898
rect 230620 204454 230940 204486
rect 230620 204218 230662 204454
rect 230898 204218 230940 204454
rect 230620 204134 230940 204218
rect 230620 203898 230662 204134
rect 230898 203898 230940 204134
rect 230620 203866 230940 203898
rect 238462 204454 238782 204486
rect 238462 204218 238504 204454
rect 238740 204218 238782 204454
rect 238462 204134 238782 204218
rect 238462 203898 238504 204134
rect 238740 203898 238782 204134
rect 238462 203866 238782 203898
rect 246304 204454 246624 204486
rect 246304 204218 246346 204454
rect 246582 204218 246624 204454
rect 246304 204134 246624 204218
rect 246304 203898 246346 204134
rect 246582 203898 246624 204134
rect 246304 203866 246624 203898
rect 256910 204454 257230 204486
rect 256910 204218 256952 204454
rect 257188 204218 257230 204454
rect 256910 204134 257230 204218
rect 256910 203898 256952 204134
rect 257188 203898 257230 204134
rect 256910 203866 257230 203898
rect 264752 204454 265072 204486
rect 264752 204218 264794 204454
rect 265030 204218 265072 204454
rect 264752 204134 265072 204218
rect 264752 203898 264794 204134
rect 265030 203898 265072 204134
rect 264752 203866 265072 203898
rect 272594 204454 272914 204486
rect 272594 204218 272636 204454
rect 272872 204218 272914 204454
rect 272594 204134 272914 204218
rect 272594 203898 272636 204134
rect 272872 203898 272914 204134
rect 272594 203866 272914 203898
rect 280436 204454 280756 204486
rect 280436 204218 280478 204454
rect 280714 204218 280756 204454
rect 280436 204134 280756 204218
rect 280436 203898 280478 204134
rect 280714 203898 280756 204134
rect 280436 203866 280756 203898
rect 184725 198174 185045 198206
rect 184725 197938 184767 198174
rect 185003 197938 185045 198174
rect 184725 197854 185045 197938
rect 184725 197618 184767 197854
rect 185003 197618 185045 197854
rect 184725 197586 185045 197618
rect 192567 198174 192887 198206
rect 192567 197938 192609 198174
rect 192845 197938 192887 198174
rect 192567 197854 192887 197938
rect 192567 197618 192609 197854
rect 192845 197618 192887 197854
rect 192567 197586 192887 197618
rect 200409 198174 200729 198206
rect 200409 197938 200451 198174
rect 200687 197938 200729 198174
rect 200409 197854 200729 197938
rect 200409 197618 200451 197854
rect 200687 197618 200729 197854
rect 200409 197586 200729 197618
rect 208251 198174 208571 198206
rect 208251 197938 208293 198174
rect 208529 197938 208571 198174
rect 208251 197854 208571 197938
rect 208251 197618 208293 197854
rect 208529 197618 208571 197854
rect 208251 197586 208571 197618
rect 218857 198174 219177 198206
rect 218857 197938 218899 198174
rect 219135 197938 219177 198174
rect 218857 197854 219177 197938
rect 218857 197618 218899 197854
rect 219135 197618 219177 197854
rect 218857 197586 219177 197618
rect 226699 198174 227019 198206
rect 226699 197938 226741 198174
rect 226977 197938 227019 198174
rect 226699 197854 227019 197938
rect 226699 197618 226741 197854
rect 226977 197618 227019 197854
rect 226699 197586 227019 197618
rect 234541 198174 234861 198206
rect 234541 197938 234583 198174
rect 234819 197938 234861 198174
rect 234541 197854 234861 197938
rect 234541 197618 234583 197854
rect 234819 197618 234861 197854
rect 234541 197586 234861 197618
rect 242383 198174 242703 198206
rect 242383 197938 242425 198174
rect 242661 197938 242703 198174
rect 242383 197854 242703 197938
rect 242383 197618 242425 197854
rect 242661 197618 242703 197854
rect 242383 197586 242703 197618
rect 252989 198174 253309 198206
rect 252989 197938 253031 198174
rect 253267 197938 253309 198174
rect 252989 197854 253309 197938
rect 252989 197618 253031 197854
rect 253267 197618 253309 197854
rect 252989 197586 253309 197618
rect 260831 198174 261151 198206
rect 260831 197938 260873 198174
rect 261109 197938 261151 198174
rect 260831 197854 261151 197938
rect 260831 197618 260873 197854
rect 261109 197618 261151 197854
rect 260831 197586 261151 197618
rect 268673 198174 268993 198206
rect 268673 197938 268715 198174
rect 268951 197938 268993 198174
rect 268673 197854 268993 197938
rect 268673 197618 268715 197854
rect 268951 197618 268993 197854
rect 268673 197586 268993 197618
rect 276515 198174 276835 198206
rect 276515 197938 276557 198174
rect 276793 197938 276835 198174
rect 276515 197854 276835 197938
rect 276515 197618 276557 197854
rect 276793 197618 276835 197854
rect 276515 197586 276835 197618
rect 188646 194454 188966 194486
rect 188646 194218 188688 194454
rect 188924 194218 188966 194454
rect 188646 194134 188966 194218
rect 188646 193898 188688 194134
rect 188924 193898 188966 194134
rect 188646 193866 188966 193898
rect 196488 194454 196808 194486
rect 196488 194218 196530 194454
rect 196766 194218 196808 194454
rect 196488 194134 196808 194218
rect 196488 193898 196530 194134
rect 196766 193898 196808 194134
rect 196488 193866 196808 193898
rect 204330 194454 204650 194486
rect 204330 194218 204372 194454
rect 204608 194218 204650 194454
rect 204330 194134 204650 194218
rect 204330 193898 204372 194134
rect 204608 193898 204650 194134
rect 204330 193866 204650 193898
rect 212172 194454 212492 194486
rect 212172 194218 212214 194454
rect 212450 194218 212492 194454
rect 212172 194134 212492 194218
rect 212172 193898 212214 194134
rect 212450 193898 212492 194134
rect 212172 193866 212492 193898
rect 222778 194454 223098 194486
rect 222778 194218 222820 194454
rect 223056 194218 223098 194454
rect 222778 194134 223098 194218
rect 222778 193898 222820 194134
rect 223056 193898 223098 194134
rect 222778 193866 223098 193898
rect 230620 194454 230940 194486
rect 230620 194218 230662 194454
rect 230898 194218 230940 194454
rect 230620 194134 230940 194218
rect 230620 193898 230662 194134
rect 230898 193898 230940 194134
rect 230620 193866 230940 193898
rect 238462 194454 238782 194486
rect 238462 194218 238504 194454
rect 238740 194218 238782 194454
rect 238462 194134 238782 194218
rect 238462 193898 238504 194134
rect 238740 193898 238782 194134
rect 238462 193866 238782 193898
rect 246304 194454 246624 194486
rect 246304 194218 246346 194454
rect 246582 194218 246624 194454
rect 246304 194134 246624 194218
rect 246304 193898 246346 194134
rect 246582 193898 246624 194134
rect 246304 193866 246624 193898
rect 256910 194454 257230 194486
rect 256910 194218 256952 194454
rect 257188 194218 257230 194454
rect 256910 194134 257230 194218
rect 256910 193898 256952 194134
rect 257188 193898 257230 194134
rect 256910 193866 257230 193898
rect 264752 194454 265072 194486
rect 264752 194218 264794 194454
rect 265030 194218 265072 194454
rect 264752 194134 265072 194218
rect 264752 193898 264794 194134
rect 265030 193898 265072 194134
rect 264752 193866 265072 193898
rect 272594 194454 272914 194486
rect 272594 194218 272636 194454
rect 272872 194218 272914 194454
rect 272594 194134 272914 194218
rect 272594 193898 272636 194134
rect 272872 193898 272914 194134
rect 272594 193866 272914 193898
rect 280436 194454 280756 194486
rect 280436 194218 280478 194454
rect 280714 194218 280756 194454
rect 280436 194134 280756 194218
rect 280436 193898 280478 194134
rect 280714 193898 280756 194134
rect 280436 193866 280756 193898
rect 281030 193221 281090 619107
rect 281947 281076 282013 281077
rect 281947 281012 281948 281076
rect 282012 281012 282013 281076
rect 281947 281011 282013 281012
rect 281763 214572 281829 214573
rect 281763 214508 281764 214572
rect 281828 214508 281829 214572
rect 281763 214507 281829 214508
rect 281027 193220 281093 193221
rect 281027 193156 281028 193220
rect 281092 193156 281093 193220
rect 281027 193155 281093 193156
rect 181394 190400 181454 191420
rect 182130 190400 182190 191420
rect 182866 190400 182926 191080
rect 183602 190400 183662 191420
rect 184338 190400 184398 191080
rect 185074 190400 185134 191080
rect 185810 190400 185870 191080
rect 186546 190400 186606 191080
rect 187282 190400 187342 191080
rect 188018 190400 188078 191080
rect 188754 190400 188814 191080
rect 189490 190400 189550 191080
rect 190226 190400 190286 191080
rect 190962 190400 191022 191080
rect 191698 190400 191758 191080
rect 192434 190400 192494 191080
rect 193170 190400 193230 191080
rect 193906 190400 193966 191080
rect 194642 190400 194702 191080
rect 195378 190400 195438 191080
rect 196114 190400 196174 191080
rect 196850 190400 196910 191080
rect 197586 190400 197646 191080
rect 198322 190400 198382 191420
rect 199058 190400 199118 191044
rect 199794 190400 199854 191044
rect 200530 190400 200590 191044
rect 201266 190400 201326 191044
rect 202002 190400 202062 191044
rect 202738 190400 202798 191044
rect 203474 190400 203534 191044
rect 204210 190400 204270 191044
rect 204946 190400 205006 191044
rect 205682 190400 205742 191044
rect 206418 190400 206478 191044
rect 207154 190400 207214 191080
rect 207890 190400 207950 191080
rect 208626 190400 208686 191080
rect 209362 190400 209422 191080
rect 210098 190770 210158 191420
rect 210098 190710 210250 190770
rect 210190 190470 210250 190710
rect 210098 190410 210250 190470
rect 210098 190400 210158 190410
rect 210834 190400 210894 191080
rect 211570 190400 211630 191080
rect 212306 190400 212366 191044
rect 215526 190400 215586 191420
rect 216262 190770 216322 191420
rect 216078 190710 216322 190770
rect 216078 190470 216138 190710
rect 216078 190410 216322 190470
rect 216262 190400 216322 190410
rect 216998 190400 217058 191420
rect 217734 190400 217794 191420
rect 218470 190400 218530 191420
rect 219206 190400 219266 191080
rect 219942 190400 220002 191420
rect 220678 190400 220738 191420
rect 221414 190400 221474 191080
rect 222150 190400 222210 191420
rect 222886 190400 222946 191080
rect 223622 190400 223682 191080
rect 224358 190400 224418 191420
rect 225094 190400 225154 191420
rect 225830 190400 225890 191420
rect 226566 190400 226626 191080
rect 227302 190400 227362 191420
rect 228038 190400 228098 191420
rect 228774 190400 228834 191080
rect 229510 190400 229570 191420
rect 230246 190400 230306 191420
rect 230982 190400 231042 191080
rect 231718 190400 231778 191420
rect 232454 190400 232514 191420
rect 233190 190400 233250 191080
rect 233926 190060 233986 191420
rect 234662 190060 234722 191080
rect 235398 190060 235458 191420
rect 236134 190060 236194 191420
rect 236870 190400 236930 191420
rect 237606 190400 237666 191420
rect 238342 190060 238402 191420
rect 239078 190400 239138 191420
rect 239814 190060 239874 191420
rect 240550 190060 240610 191420
rect 241286 190400 241346 191420
rect 242022 190060 242082 191420
rect 242758 190400 242818 191080
rect 243494 190060 243554 191420
rect 244230 190060 244290 191420
rect 244966 190400 245026 191420
rect 245702 190400 245762 191080
rect 246438 190060 246498 191044
rect 249658 190400 249718 191080
rect 250394 190400 250454 191080
rect 251130 190400 251190 191080
rect 251866 190400 251926 191080
rect 252602 190400 252662 191080
rect 253338 190400 253398 191080
rect 254074 190400 254134 191080
rect 254810 190400 254870 191080
rect 255546 190400 255606 191080
rect 256282 190400 256342 191080
rect 257018 190400 257078 191080
rect 257754 190400 257814 191080
rect 258490 190400 258550 191080
rect 259226 190400 259286 191080
rect 259962 190400 260022 191080
rect 260698 190400 260758 191080
rect 261434 190400 261494 191080
rect 262170 190400 262230 191080
rect 262906 190400 262966 191080
rect 263642 190400 263702 191080
rect 264378 190400 264438 191080
rect 265114 190400 265174 191080
rect 265850 190400 265910 191080
rect 266586 190400 266646 191080
rect 267322 190400 267382 191044
rect 268058 190400 268118 191044
rect 268794 190400 268854 191044
rect 269530 190400 269590 191044
rect 270266 190400 270326 191044
rect 271002 190400 271062 191044
rect 271738 190400 271798 191044
rect 272474 190400 272534 191044
rect 273210 190400 273270 191044
rect 273946 190400 274006 191044
rect 274682 190400 274742 191044
rect 275418 190400 275478 191044
rect 276154 190400 276214 191044
rect 276890 190400 276950 191044
rect 277626 190400 277686 191044
rect 278362 190400 278422 191044
rect 279098 190400 279158 191080
rect 279834 190400 279894 191080
rect 280570 190400 280630 191044
rect 281395 190636 281461 190637
rect 281395 190572 281396 190636
rect 281460 190572 281461 190636
rect 281395 190571 281461 190572
rect 43942 188174 44262 188206
rect 43942 187938 43984 188174
rect 44220 187938 44262 188174
rect 43942 187854 44262 187938
rect 43942 187618 43984 187854
rect 44220 187618 44262 187854
rect 43942 187586 44262 187618
rect 111539 188174 111859 188206
rect 111539 187938 111581 188174
rect 111817 187938 111859 188174
rect 111539 187854 111859 187938
rect 111539 187618 111581 187854
rect 111817 187618 111859 187854
rect 111539 187586 111859 187618
rect 179136 188174 179456 188206
rect 179136 187938 179178 188174
rect 179414 187938 179456 188174
rect 179136 187854 179456 187938
rect 179136 187618 179178 187854
rect 179414 187618 179456 187854
rect 179136 187586 179456 187618
rect 246733 188174 247053 188206
rect 246733 187938 246775 188174
rect 247011 187938 247053 188174
rect 246733 187854 247053 187938
rect 246733 187618 246775 187854
rect 247011 187618 247053 187854
rect 246733 187586 247053 187618
rect 281398 187373 281458 190571
rect 281395 187372 281461 187373
rect 281395 187308 281396 187372
rect 281460 187308 281461 187372
rect 281395 187307 281461 187308
rect 77740 184454 78060 184486
rect 77740 184218 77782 184454
rect 78018 184218 78060 184454
rect 77740 184134 78060 184218
rect 77740 183898 77782 184134
rect 78018 183898 78060 184134
rect 77740 183866 78060 183898
rect 145337 184454 145657 184486
rect 145337 184218 145379 184454
rect 145615 184218 145657 184454
rect 145337 184134 145657 184218
rect 145337 183898 145379 184134
rect 145615 183898 145657 184134
rect 145337 183866 145657 183898
rect 212934 184454 213254 184486
rect 212934 184218 212976 184454
rect 213212 184218 213254 184454
rect 212934 184134 213254 184218
rect 212934 183898 212976 184134
rect 213212 183898 213254 184134
rect 212934 183866 213254 183898
rect 280531 184454 280851 184486
rect 280531 184218 280573 184454
rect 280809 184218 280851 184454
rect 280531 184134 280851 184218
rect 280531 183898 280573 184134
rect 280809 183898 280851 184134
rect 280531 183866 280851 183898
rect 281027 182476 281093 182477
rect 281027 182412 281028 182476
rect 281092 182412 281093 182476
rect 281027 182411 281093 182412
rect 10734 134758 10794 179520
rect 11470 134758 11530 179520
rect 12206 134758 12266 179520
rect 12942 134690 13002 179520
rect 13678 134690 13738 179520
rect 14414 134758 14474 179520
rect 15150 134758 15210 179520
rect 15886 134690 15946 179520
rect 16622 134300 16682 179520
rect 17358 134300 17418 179520
rect 18094 134300 18154 179520
rect 18830 134300 18890 179520
rect 19566 134300 19626 179520
rect 20302 134300 20362 179520
rect 21038 134300 21098 179520
rect 21774 134300 21834 179520
rect 22510 134758 22570 179520
rect 23246 134758 23306 179520
rect 23982 134758 24042 179520
rect 24718 134300 24778 179520
rect 25454 134758 25514 179520
rect 26190 179210 26250 179520
rect 26006 179150 26250 179210
rect 26006 135690 26066 179150
rect 26006 135630 26250 135690
rect 26190 134758 26250 135630
rect 26926 134640 26986 179520
rect 27662 134300 27722 179520
rect 28398 134758 28458 179860
rect 29134 134640 29194 179520
rect 29870 134640 29930 179520
rect 30606 134758 30666 179520
rect 31342 134758 31402 179520
rect 32078 134690 32138 179860
rect 32814 134640 32874 179520
rect 33550 134640 33610 179520
rect 34286 134812 34346 179860
rect 35022 134640 35082 179520
rect 35758 134640 35818 179520
rect 36494 134640 36554 179860
rect 37230 134640 37290 179520
rect 37966 134640 38026 179520
rect 38702 134640 38762 179520
rect 39438 134640 39498 179520
rect 40174 134690 40234 179520
rect 40910 134795 40970 179520
rect 41646 134812 41706 179520
rect 44866 178840 44926 179520
rect 45602 178840 45662 179520
rect 46338 178840 46398 179520
rect 47074 178840 47134 179520
rect 47810 178840 47870 179520
rect 48546 178840 48606 179520
rect 49282 178840 49342 179520
rect 50018 178840 50078 179520
rect 50754 178840 50814 179520
rect 51490 178840 51550 179520
rect 52226 178840 52286 179520
rect 52962 178840 53022 179520
rect 53698 178840 53758 179520
rect 54434 178840 54494 179520
rect 55170 178840 55230 179520
rect 55906 178840 55966 179520
rect 56642 178840 56702 179520
rect 57378 178840 57438 179520
rect 58114 178840 58174 179520
rect 58850 178840 58910 179520
rect 59586 178840 59646 179520
rect 60322 178840 60382 179520
rect 61058 178840 61118 179520
rect 61794 178840 61854 179520
rect 62530 178876 62590 179520
rect 63266 178876 63326 179520
rect 64002 178876 64062 179520
rect 64738 178876 64798 179520
rect 65474 178876 65534 179520
rect 66210 178876 66270 179520
rect 66946 178876 67006 179520
rect 67682 178876 67742 179520
rect 68418 178876 68478 179520
rect 69154 178876 69214 179520
rect 69890 178876 69950 179520
rect 70626 178876 70686 179520
rect 71362 178840 71422 179520
rect 72098 178840 72158 179520
rect 72834 178840 72894 179520
rect 73570 178840 73630 179520
rect 74306 178840 74366 179520
rect 75042 178500 75102 179520
rect 75778 178876 75838 179520
rect 78998 178840 79058 179520
rect 79734 178840 79794 179520
rect 80470 178840 80530 179520
rect 81206 178840 81266 179520
rect 81942 178840 82002 179520
rect 82678 178840 82738 179520
rect 83414 178840 83474 179520
rect 84150 178840 84210 179520
rect 84886 178840 84946 179520
rect 85622 178840 85682 179520
rect 86358 178840 86418 179520
rect 87094 178840 87154 179520
rect 87830 178840 87890 179520
rect 88566 178840 88626 179520
rect 89302 178840 89362 179520
rect 90038 178840 90098 179520
rect 90774 178840 90834 179520
rect 91510 178840 91570 179520
rect 92246 178840 92306 179520
rect 92982 178840 93042 179520
rect 93718 178840 93778 179520
rect 94454 178840 94514 179520
rect 95190 178840 95250 179520
rect 95926 178840 95986 179520
rect 96662 178876 96722 179520
rect 97398 178876 97458 179520
rect 98134 178876 98194 179520
rect 98870 178876 98930 179520
rect 99606 178876 99666 179520
rect 100342 178876 100402 179520
rect 101078 178876 101138 179520
rect 101814 178876 101874 179520
rect 102550 178876 102610 179520
rect 103286 178876 103346 179860
rect 104022 178840 104082 179520
rect 104758 178840 104818 179860
rect 105494 178840 105554 179520
rect 106230 178840 106290 179860
rect 106966 178876 107026 179860
rect 107702 178876 107762 179520
rect 108438 178840 108498 179520
rect 109174 178500 109234 179520
rect 109910 178876 109970 179860
rect 113130 178840 113190 179520
rect 113866 178840 113926 179520
rect 114602 178840 114662 179520
rect 115338 178840 115398 179520
rect 116074 178840 116134 179520
rect 116810 178840 116870 179520
rect 117546 178840 117606 179520
rect 118282 178840 118342 179520
rect 119018 178840 119078 179520
rect 119754 178840 119814 179520
rect 120490 178840 120550 179520
rect 121226 178840 121286 179520
rect 121962 178840 122022 179520
rect 122698 178840 122758 179520
rect 123434 178840 123494 179520
rect 124170 178840 124230 179520
rect 124906 178840 124966 179520
rect 125642 178500 125702 179520
rect 126378 178840 126438 179520
rect 127114 178500 127174 179520
rect 127850 178840 127910 179520
rect 128586 178840 128646 179520
rect 129322 178500 129382 179520
rect 130058 178500 130118 179520
rect 130794 178840 130854 179520
rect 131530 178876 131590 179520
rect 132266 178840 132326 179520
rect 133002 178840 133062 179520
rect 133738 178840 133798 179520
rect 134474 178840 134534 179520
rect 135210 178840 135270 179520
rect 135946 178840 136006 179520
rect 136682 178840 136742 179520
rect 137418 178840 137478 179520
rect 138154 178840 138214 179520
rect 138890 178840 138950 179520
rect 139626 178840 139686 179520
rect 140362 178840 140422 179520
rect 141098 178840 141158 179520
rect 141834 178840 141894 179520
rect 142570 178840 142630 179520
rect 143306 178876 143366 179520
rect 144042 178876 144102 179520
rect 147262 178840 147322 179520
rect 147998 178840 148058 179520
rect 148734 178840 148794 179520
rect 149470 178840 149530 179860
rect 150206 178840 150266 179520
rect 150942 178840 151002 179520
rect 151678 178840 151738 179520
rect 152414 178840 152474 179520
rect 153150 178840 153210 179520
rect 153886 178840 153946 179860
rect 154622 178840 154682 179860
rect 155358 178840 155418 179520
rect 156094 178840 156154 179520
rect 156830 178840 156890 179520
rect 157566 178840 157626 179520
rect 158302 178840 158362 179860
rect 159038 178500 159098 179520
rect 159774 178500 159834 179520
rect 160510 178500 160570 179520
rect 161246 178500 161306 179520
rect 161982 178500 162042 179520
rect 162718 178500 162778 179860
rect 163454 178500 163514 179860
rect 164190 178500 164250 179860
rect 164926 178840 164986 179520
rect 165662 178840 165722 179860
rect 166398 178840 166458 179520
rect 167134 178840 167194 179520
rect 167870 178840 167930 179520
rect 168606 178840 168666 179520
rect 169342 178840 169402 179520
rect 170078 178840 170138 179520
rect 170814 178840 170874 179520
rect 171550 178840 171610 179520
rect 172286 178840 172346 179520
rect 173022 178840 173082 179520
rect 173758 178840 173818 179520
rect 174494 178840 174554 179520
rect 175230 178840 175290 179520
rect 175966 178840 176026 179520
rect 176702 178840 176762 179520
rect 177438 178500 177498 179520
rect 178174 178876 178234 179520
rect 180658 179346 180718 179520
rect 181394 179346 181454 179520
rect 182130 179349 182190 179520
rect 182866 179349 182926 179520
rect 183602 179349 183662 179520
rect 184338 179349 184398 179520
rect 185074 179349 185134 179520
rect 182127 179348 182193 179349
rect 182127 179346 182128 179348
rect 180658 179286 182128 179346
rect 182127 179284 182128 179286
rect 182192 179284 182193 179348
rect 182127 179283 182193 179284
rect 182863 179348 182929 179349
rect 182863 179284 182864 179348
rect 182928 179284 182929 179348
rect 182863 179283 182929 179284
rect 183599 179348 183665 179349
rect 183599 179284 183600 179348
rect 183664 179284 183665 179348
rect 183599 179283 183665 179284
rect 184335 179348 184401 179349
rect 184335 179284 184336 179348
rect 184400 179284 184401 179348
rect 184335 179283 184401 179284
rect 185071 179348 185137 179349
rect 185071 179284 185072 179348
rect 185136 179284 185137 179348
rect 185071 179283 185137 179284
rect 185810 179213 185870 179520
rect 186546 179349 186606 179520
rect 187282 179349 187342 179520
rect 188018 179349 188078 179520
rect 188754 179349 188814 179520
rect 189490 179349 189550 179520
rect 190226 179349 190286 179520
rect 186543 179348 186609 179349
rect 186543 179284 186544 179348
rect 186608 179284 186609 179348
rect 186543 179283 186609 179284
rect 187279 179348 187345 179349
rect 187279 179284 187280 179348
rect 187344 179284 187345 179348
rect 187279 179283 187345 179284
rect 188015 179348 188081 179349
rect 188015 179284 188016 179348
rect 188080 179284 188081 179348
rect 188015 179283 188081 179284
rect 188751 179348 188817 179349
rect 188751 179284 188752 179348
rect 188816 179284 188817 179348
rect 188751 179283 188817 179284
rect 189487 179348 189553 179349
rect 189487 179284 189488 179348
rect 189552 179284 189553 179348
rect 189487 179283 189553 179284
rect 190223 179348 190289 179349
rect 190223 179284 190224 179348
rect 190288 179284 190289 179348
rect 190223 179283 190289 179284
rect 190962 179213 191022 179520
rect 191698 179349 191758 179520
rect 192434 179349 192494 179520
rect 193170 179349 193230 179520
rect 193906 179349 193966 179520
rect 194642 179349 194702 179520
rect 195378 179349 195438 179520
rect 196114 179349 196174 179520
rect 196850 179349 196910 179520
rect 197586 179349 197646 179520
rect 198322 179349 198382 179520
rect 214790 179349 214850 179520
rect 215526 179349 215586 179520
rect 216262 179349 216322 179520
rect 216998 179349 217058 179520
rect 217734 179349 217794 179520
rect 218470 179349 218530 179520
rect 219206 179349 219266 179520
rect 219942 179349 220002 179860
rect 220678 179550 220738 179860
rect 220678 179490 220922 179550
rect 220862 179349 220922 179490
rect 221414 179349 221474 179860
rect 224358 179550 224418 179860
rect 225830 179550 225890 179860
rect 226566 179550 226626 179860
rect 228038 179550 228098 179860
rect 230246 179550 230306 179860
rect 232454 179550 232514 179860
rect 222150 179349 222210 179520
rect 222886 179349 222946 179520
rect 223622 179349 223682 179520
rect 223806 179490 224970 179550
rect 191695 179348 191761 179349
rect 191695 179284 191696 179348
rect 191760 179284 191761 179348
rect 191695 179283 191761 179284
rect 192431 179348 192497 179349
rect 192431 179284 192432 179348
rect 192496 179284 192497 179348
rect 192431 179283 192497 179284
rect 193167 179348 193233 179349
rect 193167 179284 193168 179348
rect 193232 179284 193233 179348
rect 193167 179283 193233 179284
rect 193903 179348 193969 179349
rect 193903 179284 193904 179348
rect 193968 179284 193969 179348
rect 193903 179283 193969 179284
rect 194639 179348 194705 179349
rect 194639 179284 194640 179348
rect 194704 179284 194705 179348
rect 194639 179283 194705 179284
rect 195375 179348 195441 179349
rect 195375 179284 195376 179348
rect 195440 179284 195441 179348
rect 195375 179283 195441 179284
rect 196111 179348 196177 179349
rect 196111 179284 196112 179348
rect 196176 179284 196177 179348
rect 196111 179283 196177 179284
rect 196847 179348 196913 179349
rect 196847 179284 196848 179348
rect 196912 179284 196913 179348
rect 196847 179283 196913 179284
rect 197583 179348 197649 179349
rect 197583 179284 197584 179348
rect 197648 179284 197649 179348
rect 197583 179283 197649 179284
rect 198319 179348 198385 179349
rect 198319 179284 198320 179348
rect 198384 179284 198385 179348
rect 198319 179283 198385 179284
rect 214787 179348 214853 179349
rect 214787 179284 214788 179348
rect 214852 179284 214853 179348
rect 214787 179283 214853 179284
rect 215523 179348 215589 179349
rect 215523 179284 215524 179348
rect 215588 179284 215589 179348
rect 215523 179283 215589 179284
rect 216259 179348 216325 179349
rect 216259 179284 216260 179348
rect 216324 179284 216325 179348
rect 216259 179283 216325 179284
rect 216995 179348 217061 179349
rect 216995 179284 216996 179348
rect 217060 179284 217061 179348
rect 216995 179283 217061 179284
rect 217731 179348 217797 179349
rect 217731 179284 217732 179348
rect 217796 179284 217797 179348
rect 217731 179283 217797 179284
rect 218467 179348 218533 179349
rect 218467 179284 218468 179348
rect 218532 179284 218533 179348
rect 218467 179283 218533 179284
rect 219203 179348 219269 179349
rect 219203 179284 219204 179348
rect 219268 179284 219269 179348
rect 219203 179283 219269 179284
rect 219939 179348 220005 179349
rect 219939 179284 219940 179348
rect 220004 179284 220005 179348
rect 219939 179283 220005 179284
rect 220859 179348 220925 179349
rect 220859 179284 220860 179348
rect 220924 179284 220925 179348
rect 220859 179283 220925 179284
rect 221411 179348 221477 179349
rect 221411 179284 221412 179348
rect 221476 179284 221477 179348
rect 221411 179283 221477 179284
rect 222147 179348 222213 179349
rect 222147 179284 222148 179348
rect 222212 179284 222213 179348
rect 222147 179283 222213 179284
rect 222883 179348 222949 179349
rect 222883 179284 222884 179348
rect 222948 179284 222949 179348
rect 222883 179283 222949 179284
rect 223619 179348 223685 179349
rect 223619 179284 223620 179348
rect 223684 179346 223685 179348
rect 223806 179346 223866 179490
rect 223684 179286 223866 179346
rect 224910 179346 224970 179490
rect 225094 179346 225154 179520
rect 225278 179490 227178 179550
rect 225278 179346 225338 179490
rect 224910 179286 225338 179346
rect 227118 179346 227178 179490
rect 227302 179346 227362 179520
rect 227486 179490 228650 179550
rect 227486 179346 227546 179490
rect 227118 179286 227546 179346
rect 228590 179346 228650 179490
rect 228774 179346 228834 179520
rect 228958 179490 229386 179550
rect 228958 179346 229018 179490
rect 228590 179286 229018 179346
rect 229326 179346 229386 179490
rect 229510 179346 229570 179520
rect 229694 179490 230858 179550
rect 229694 179346 229754 179490
rect 229326 179286 229754 179346
rect 230798 179346 230858 179490
rect 230982 179346 231042 179520
rect 231166 179490 231594 179550
rect 231166 179346 231226 179490
rect 230798 179286 231226 179346
rect 231534 179346 231594 179490
rect 231718 179346 231778 179520
rect 231902 179490 232514 179550
rect 231902 179346 231962 179490
rect 248922 179349 248982 179520
rect 249658 179349 249718 179520
rect 250394 179349 250454 179520
rect 251130 179349 251190 179520
rect 251866 179349 251926 179520
rect 252602 179349 252662 179520
rect 253338 179349 253398 179520
rect 254074 179349 254134 179520
rect 254810 179349 254870 179520
rect 255546 179349 255606 179520
rect 256282 179349 256342 179520
rect 257018 179349 257078 179520
rect 257754 179349 257814 179520
rect 258490 179349 258550 179520
rect 259226 179349 259286 179520
rect 259962 179349 260022 179520
rect 260698 179349 260758 179520
rect 261434 179349 261494 179520
rect 262170 179349 262230 179520
rect 262906 179349 262966 179520
rect 263642 179349 263702 179520
rect 264378 179349 264438 179520
rect 265114 179349 265174 179520
rect 265850 179349 265910 179520
rect 266586 179349 266646 179520
rect 231534 179286 231962 179346
rect 248919 179348 248985 179349
rect 223684 179284 223685 179286
rect 223619 179283 223685 179284
rect 248919 179284 248920 179348
rect 248984 179284 248985 179348
rect 248919 179283 248985 179284
rect 249655 179348 249721 179349
rect 249655 179284 249656 179348
rect 249720 179284 249721 179348
rect 249655 179283 249721 179284
rect 250391 179348 250457 179349
rect 250391 179284 250392 179348
rect 250456 179284 250457 179348
rect 250391 179283 250457 179284
rect 251127 179348 251193 179349
rect 251127 179284 251128 179348
rect 251192 179284 251193 179348
rect 251127 179283 251193 179284
rect 251863 179348 251929 179349
rect 251863 179284 251864 179348
rect 251928 179284 251929 179348
rect 251863 179283 251929 179284
rect 252599 179348 252665 179349
rect 252599 179284 252600 179348
rect 252664 179284 252665 179348
rect 252599 179283 252665 179284
rect 253335 179348 253401 179349
rect 253335 179284 253336 179348
rect 253400 179284 253401 179348
rect 253335 179283 253401 179284
rect 254071 179348 254137 179349
rect 254071 179284 254072 179348
rect 254136 179284 254137 179348
rect 254071 179283 254137 179284
rect 254807 179348 254873 179349
rect 254807 179284 254808 179348
rect 254872 179284 254873 179348
rect 254807 179283 254873 179284
rect 255543 179348 255609 179349
rect 255543 179284 255544 179348
rect 255608 179284 255609 179348
rect 255543 179283 255609 179284
rect 256279 179348 256345 179349
rect 256279 179284 256280 179348
rect 256344 179284 256345 179348
rect 256279 179283 256345 179284
rect 257015 179348 257081 179349
rect 257015 179284 257016 179348
rect 257080 179284 257081 179348
rect 257015 179283 257081 179284
rect 257751 179348 257817 179349
rect 257751 179284 257752 179348
rect 257816 179284 257817 179348
rect 257751 179283 257817 179284
rect 258487 179348 258553 179349
rect 258487 179284 258488 179348
rect 258552 179284 258553 179348
rect 258487 179283 258553 179284
rect 259223 179348 259289 179349
rect 259223 179284 259224 179348
rect 259288 179284 259289 179348
rect 259223 179283 259289 179284
rect 259959 179348 260025 179349
rect 259959 179284 259960 179348
rect 260024 179284 260025 179348
rect 259959 179283 260025 179284
rect 260695 179348 260761 179349
rect 260695 179284 260696 179348
rect 260760 179284 260761 179348
rect 260695 179283 260761 179284
rect 261431 179348 261497 179349
rect 261431 179284 261432 179348
rect 261496 179284 261497 179348
rect 261431 179283 261497 179284
rect 262167 179348 262233 179349
rect 262167 179284 262168 179348
rect 262232 179284 262233 179348
rect 262167 179283 262233 179284
rect 262903 179348 262969 179349
rect 262903 179284 262904 179348
rect 262968 179284 262969 179348
rect 262903 179283 262969 179284
rect 263639 179348 263705 179349
rect 263639 179284 263640 179348
rect 263704 179284 263705 179348
rect 263639 179283 263705 179284
rect 264375 179348 264441 179349
rect 264375 179284 264376 179348
rect 264440 179284 264441 179348
rect 264375 179283 264441 179284
rect 265111 179348 265177 179349
rect 265111 179284 265112 179348
rect 265176 179284 265177 179348
rect 265111 179283 265177 179284
rect 265847 179348 265913 179349
rect 265847 179284 265848 179348
rect 265912 179284 265913 179348
rect 265847 179283 265913 179284
rect 266583 179348 266649 179349
rect 266583 179284 266584 179348
rect 266648 179284 266649 179348
rect 266583 179283 266649 179284
rect 185807 179212 185873 179213
rect 185807 179148 185808 179212
rect 185872 179148 185873 179212
rect 185807 179147 185873 179148
rect 190959 179212 191025 179213
rect 190959 179148 190960 179212
rect 191024 179148 191025 179212
rect 190959 179147 191025 179148
rect 279003 179212 279069 179213
rect 279003 179148 279004 179212
rect 279068 179148 279069 179212
rect 279003 179147 279069 179148
rect 48197 177879 48517 177936
rect 48197 177643 48239 177879
rect 48475 177643 48517 177879
rect 48197 177586 48517 177643
rect 56039 177879 56359 177936
rect 56039 177643 56081 177879
rect 56317 177643 56359 177879
rect 56039 177586 56359 177643
rect 63881 177879 64201 177936
rect 63881 177643 63923 177879
rect 64159 177643 64201 177879
rect 63881 177586 64201 177643
rect 71723 177879 72043 177936
rect 71723 177643 71765 177879
rect 72001 177643 72043 177879
rect 71723 177586 72043 177643
rect 82329 177879 82649 177936
rect 82329 177643 82371 177879
rect 82607 177643 82649 177879
rect 82329 177586 82649 177643
rect 90171 177879 90491 177936
rect 90171 177643 90213 177879
rect 90449 177643 90491 177879
rect 90171 177586 90491 177643
rect 98013 177879 98333 177936
rect 98013 177643 98055 177879
rect 98291 177643 98333 177879
rect 98013 177586 98333 177643
rect 105855 177879 106175 177936
rect 105855 177643 105897 177879
rect 106133 177643 106175 177879
rect 105855 177586 106175 177643
rect 116461 177879 116781 177936
rect 116461 177643 116503 177879
rect 116739 177643 116781 177879
rect 116461 177586 116781 177643
rect 124303 177879 124623 177936
rect 124303 177643 124345 177879
rect 124581 177643 124623 177879
rect 124303 177586 124623 177643
rect 132145 177879 132465 177936
rect 132145 177643 132187 177879
rect 132423 177643 132465 177879
rect 132145 177586 132465 177643
rect 139987 177879 140307 177936
rect 139987 177643 140029 177879
rect 140265 177643 140307 177879
rect 139987 177586 140307 177643
rect 149936 177879 150256 177936
rect 149936 177643 149978 177879
rect 150214 177643 150256 177879
rect 149936 177586 150256 177643
rect 180656 177879 180976 177936
rect 180656 177643 180698 177879
rect 180934 177643 180976 177879
rect 180656 177586 180976 177643
rect 211376 177879 211696 177936
rect 211376 177643 211418 177879
rect 211654 177643 211696 177879
rect 211376 177586 211696 177643
rect 242096 177879 242416 177936
rect 242096 177643 242138 177879
rect 242374 177643 242416 177879
rect 242096 177586 242416 177643
rect 272816 177879 273136 177936
rect 272816 177643 272858 177879
rect 273094 177643 273136 177879
rect 272816 177586 273136 177643
rect 52118 174454 52438 174486
rect 52118 174218 52160 174454
rect 52396 174218 52438 174454
rect 52118 174134 52438 174218
rect 52118 173898 52160 174134
rect 52396 173898 52438 174134
rect 52118 173866 52438 173898
rect 59960 174454 60280 174486
rect 59960 174218 60002 174454
rect 60238 174218 60280 174454
rect 59960 174134 60280 174218
rect 59960 173898 60002 174134
rect 60238 173898 60280 174134
rect 59960 173866 60280 173898
rect 67802 174454 68122 174486
rect 67802 174218 67844 174454
rect 68080 174218 68122 174454
rect 67802 174134 68122 174218
rect 67802 173898 67844 174134
rect 68080 173898 68122 174134
rect 67802 173866 68122 173898
rect 75644 174454 75964 174486
rect 75644 174218 75686 174454
rect 75922 174218 75964 174454
rect 75644 174134 75964 174218
rect 75644 173898 75686 174134
rect 75922 173898 75964 174134
rect 75644 173866 75964 173898
rect 86250 174454 86570 174486
rect 86250 174218 86292 174454
rect 86528 174218 86570 174454
rect 86250 174134 86570 174218
rect 86250 173898 86292 174134
rect 86528 173898 86570 174134
rect 86250 173866 86570 173898
rect 94092 174454 94412 174486
rect 94092 174218 94134 174454
rect 94370 174218 94412 174454
rect 94092 174134 94412 174218
rect 94092 173898 94134 174134
rect 94370 173898 94412 174134
rect 94092 173866 94412 173898
rect 101934 174454 102254 174486
rect 101934 174218 101976 174454
rect 102212 174218 102254 174454
rect 101934 174134 102254 174218
rect 101934 173898 101976 174134
rect 102212 173898 102254 174134
rect 101934 173866 102254 173898
rect 109776 174454 110096 174486
rect 109776 174218 109818 174454
rect 110054 174218 110096 174454
rect 109776 174134 110096 174218
rect 109776 173898 109818 174134
rect 110054 173898 110096 174134
rect 109776 173866 110096 173898
rect 120382 174454 120702 174486
rect 120382 174218 120424 174454
rect 120660 174218 120702 174454
rect 120382 174134 120702 174218
rect 120382 173898 120424 174134
rect 120660 173898 120702 174134
rect 120382 173866 120702 173898
rect 128224 174454 128544 174486
rect 128224 174218 128266 174454
rect 128502 174218 128544 174454
rect 128224 174134 128544 174218
rect 128224 173898 128266 174134
rect 128502 173898 128544 174134
rect 128224 173866 128544 173898
rect 136066 174454 136386 174486
rect 136066 174218 136108 174454
rect 136344 174218 136386 174454
rect 136066 174134 136386 174218
rect 136066 173898 136108 174134
rect 136344 173898 136386 174134
rect 136066 173866 136386 173898
rect 143908 174454 144228 174486
rect 143908 174218 143950 174454
rect 144186 174218 144228 174454
rect 143908 174134 144228 174218
rect 143908 173898 143950 174134
rect 144186 173898 144228 174134
rect 143908 173866 144228 173898
rect 165296 174454 165616 174486
rect 165296 174218 165338 174454
rect 165574 174218 165616 174454
rect 165296 174134 165616 174218
rect 165296 173898 165338 174134
rect 165574 173898 165616 174134
rect 165296 173866 165616 173898
rect 196016 174454 196336 174486
rect 196016 174218 196058 174454
rect 196294 174218 196336 174454
rect 196016 174134 196336 174218
rect 196016 173898 196058 174134
rect 196294 173898 196336 174134
rect 196016 173866 196336 173898
rect 226736 174454 227056 174486
rect 226736 174218 226778 174454
rect 227014 174218 227056 174454
rect 226736 174134 227056 174218
rect 226736 173898 226778 174134
rect 227014 173898 227056 174134
rect 226736 173866 227056 173898
rect 257456 174454 257776 174486
rect 257456 174218 257498 174454
rect 257734 174218 257776 174454
rect 257456 174134 257776 174218
rect 257456 173898 257498 174134
rect 257734 173898 257776 174134
rect 257456 173866 257776 173898
rect 48197 168174 48517 168206
rect 48197 167938 48239 168174
rect 48475 167938 48517 168174
rect 48197 167854 48517 167938
rect 48197 167618 48239 167854
rect 48475 167618 48517 167854
rect 48197 167586 48517 167618
rect 56039 168174 56359 168206
rect 56039 167938 56081 168174
rect 56317 167938 56359 168174
rect 56039 167854 56359 167938
rect 56039 167618 56081 167854
rect 56317 167618 56359 167854
rect 56039 167586 56359 167618
rect 63881 168174 64201 168206
rect 63881 167938 63923 168174
rect 64159 167938 64201 168174
rect 63881 167854 64201 167938
rect 63881 167618 63923 167854
rect 64159 167618 64201 167854
rect 63881 167586 64201 167618
rect 71723 168174 72043 168206
rect 71723 167938 71765 168174
rect 72001 167938 72043 168174
rect 71723 167854 72043 167938
rect 71723 167618 71765 167854
rect 72001 167618 72043 167854
rect 71723 167586 72043 167618
rect 82329 168174 82649 168206
rect 82329 167938 82371 168174
rect 82607 167938 82649 168174
rect 82329 167854 82649 167938
rect 82329 167618 82371 167854
rect 82607 167618 82649 167854
rect 82329 167586 82649 167618
rect 90171 168174 90491 168206
rect 90171 167938 90213 168174
rect 90449 167938 90491 168174
rect 90171 167854 90491 167938
rect 90171 167618 90213 167854
rect 90449 167618 90491 167854
rect 90171 167586 90491 167618
rect 98013 168174 98333 168206
rect 98013 167938 98055 168174
rect 98291 167938 98333 168174
rect 98013 167854 98333 167938
rect 98013 167618 98055 167854
rect 98291 167618 98333 167854
rect 98013 167586 98333 167618
rect 105855 168174 106175 168206
rect 105855 167938 105897 168174
rect 106133 167938 106175 168174
rect 105855 167854 106175 167938
rect 105855 167618 105897 167854
rect 106133 167618 106175 167854
rect 105855 167586 106175 167618
rect 116461 168174 116781 168206
rect 116461 167938 116503 168174
rect 116739 167938 116781 168174
rect 116461 167854 116781 167938
rect 116461 167618 116503 167854
rect 116739 167618 116781 167854
rect 116461 167586 116781 167618
rect 124303 168174 124623 168206
rect 124303 167938 124345 168174
rect 124581 167938 124623 168174
rect 124303 167854 124623 167938
rect 124303 167618 124345 167854
rect 124581 167618 124623 167854
rect 124303 167586 124623 167618
rect 132145 168174 132465 168206
rect 132145 167938 132187 168174
rect 132423 167938 132465 168174
rect 132145 167854 132465 167938
rect 132145 167618 132187 167854
rect 132423 167618 132465 167854
rect 132145 167586 132465 167618
rect 139987 168174 140307 168206
rect 139987 167938 140029 168174
rect 140265 167938 140307 168174
rect 139987 167854 140307 167938
rect 139987 167618 140029 167854
rect 140265 167618 140307 167854
rect 139987 167586 140307 167618
rect 149936 168174 150256 168206
rect 149936 167938 149978 168174
rect 150214 167938 150256 168174
rect 149936 167854 150256 167938
rect 149936 167618 149978 167854
rect 150214 167618 150256 167854
rect 149936 167586 150256 167618
rect 180656 168174 180976 168206
rect 180656 167938 180698 168174
rect 180934 167938 180976 168174
rect 180656 167854 180976 167938
rect 180656 167618 180698 167854
rect 180934 167618 180976 167854
rect 180656 167586 180976 167618
rect 211376 168174 211696 168206
rect 211376 167938 211418 168174
rect 211654 167938 211696 168174
rect 211376 167854 211696 167938
rect 211376 167618 211418 167854
rect 211654 167618 211696 167854
rect 211376 167586 211696 167618
rect 242096 168174 242416 168206
rect 242096 167938 242138 168174
rect 242374 167938 242416 168174
rect 242096 167854 242416 167938
rect 242096 167618 242138 167854
rect 242374 167618 242416 167854
rect 242096 167586 242416 167618
rect 272816 168174 273136 168206
rect 272816 167938 272858 168174
rect 273094 167938 273136 168174
rect 272816 167854 273136 167938
rect 272816 167618 272858 167854
rect 273094 167618 273136 167854
rect 272816 167586 273136 167618
rect 52118 164454 52438 164486
rect 52118 164218 52160 164454
rect 52396 164218 52438 164454
rect 52118 164134 52438 164218
rect 52118 163898 52160 164134
rect 52396 163898 52438 164134
rect 52118 163866 52438 163898
rect 59960 164454 60280 164486
rect 59960 164218 60002 164454
rect 60238 164218 60280 164454
rect 59960 164134 60280 164218
rect 59960 163898 60002 164134
rect 60238 163898 60280 164134
rect 59960 163866 60280 163898
rect 67802 164454 68122 164486
rect 67802 164218 67844 164454
rect 68080 164218 68122 164454
rect 67802 164134 68122 164218
rect 67802 163898 67844 164134
rect 68080 163898 68122 164134
rect 67802 163866 68122 163898
rect 75644 164454 75964 164486
rect 75644 164218 75686 164454
rect 75922 164218 75964 164454
rect 75644 164134 75964 164218
rect 75644 163898 75686 164134
rect 75922 163898 75964 164134
rect 75644 163866 75964 163898
rect 86250 164454 86570 164486
rect 86250 164218 86292 164454
rect 86528 164218 86570 164454
rect 86250 164134 86570 164218
rect 86250 163898 86292 164134
rect 86528 163898 86570 164134
rect 86250 163866 86570 163898
rect 94092 164454 94412 164486
rect 94092 164218 94134 164454
rect 94370 164218 94412 164454
rect 94092 164134 94412 164218
rect 94092 163898 94134 164134
rect 94370 163898 94412 164134
rect 94092 163866 94412 163898
rect 101934 164454 102254 164486
rect 101934 164218 101976 164454
rect 102212 164218 102254 164454
rect 101934 164134 102254 164218
rect 101934 163898 101976 164134
rect 102212 163898 102254 164134
rect 101934 163866 102254 163898
rect 109776 164454 110096 164486
rect 109776 164218 109818 164454
rect 110054 164218 110096 164454
rect 109776 164134 110096 164218
rect 109776 163898 109818 164134
rect 110054 163898 110096 164134
rect 109776 163866 110096 163898
rect 120382 164454 120702 164486
rect 120382 164218 120424 164454
rect 120660 164218 120702 164454
rect 120382 164134 120702 164218
rect 120382 163898 120424 164134
rect 120660 163898 120702 164134
rect 120382 163866 120702 163898
rect 128224 164454 128544 164486
rect 128224 164218 128266 164454
rect 128502 164218 128544 164454
rect 128224 164134 128544 164218
rect 128224 163898 128266 164134
rect 128502 163898 128544 164134
rect 128224 163866 128544 163898
rect 136066 164454 136386 164486
rect 136066 164218 136108 164454
rect 136344 164218 136386 164454
rect 136066 164134 136386 164218
rect 136066 163898 136108 164134
rect 136344 163898 136386 164134
rect 136066 163866 136386 163898
rect 143908 164454 144228 164486
rect 143908 164218 143950 164454
rect 144186 164218 144228 164454
rect 143908 164134 144228 164218
rect 143908 163898 143950 164134
rect 144186 163898 144228 164134
rect 143908 163866 144228 163898
rect 165296 164454 165616 164486
rect 165296 164218 165338 164454
rect 165574 164218 165616 164454
rect 165296 164134 165616 164218
rect 165296 163898 165338 164134
rect 165574 163898 165616 164134
rect 165296 163866 165616 163898
rect 196016 164454 196336 164486
rect 196016 164218 196058 164454
rect 196294 164218 196336 164454
rect 196016 164134 196336 164218
rect 196016 163898 196058 164134
rect 196294 163898 196336 164134
rect 196016 163866 196336 163898
rect 226736 164454 227056 164486
rect 226736 164218 226778 164454
rect 227014 164218 227056 164454
rect 226736 164134 227056 164218
rect 226736 163898 226778 164134
rect 227014 163898 227056 164134
rect 226736 163866 227056 163898
rect 257456 164454 257776 164486
rect 257456 164218 257498 164454
rect 257734 164218 257776 164454
rect 257456 164134 257776 164218
rect 257456 163898 257498 164134
rect 257734 163898 257776 164134
rect 257456 163866 257776 163898
rect 277772 164454 278092 164486
rect 277772 164218 277814 164454
rect 278050 164218 278092 164454
rect 277772 164134 278092 164218
rect 277772 163898 277814 164134
rect 278050 163898 278092 164134
rect 277772 163866 278092 163898
rect 48197 158174 48517 158206
rect 48197 157938 48239 158174
rect 48475 157938 48517 158174
rect 48197 157854 48517 157938
rect 48197 157618 48239 157854
rect 48475 157618 48517 157854
rect 48197 157586 48517 157618
rect 56039 158174 56359 158206
rect 56039 157938 56081 158174
rect 56317 157938 56359 158174
rect 56039 157854 56359 157938
rect 56039 157618 56081 157854
rect 56317 157618 56359 157854
rect 56039 157586 56359 157618
rect 63881 158174 64201 158206
rect 63881 157938 63923 158174
rect 64159 157938 64201 158174
rect 63881 157854 64201 157938
rect 63881 157618 63923 157854
rect 64159 157618 64201 157854
rect 63881 157586 64201 157618
rect 71723 158174 72043 158206
rect 71723 157938 71765 158174
rect 72001 157938 72043 158174
rect 71723 157854 72043 157938
rect 71723 157618 71765 157854
rect 72001 157618 72043 157854
rect 71723 157586 72043 157618
rect 82329 158174 82649 158206
rect 82329 157938 82371 158174
rect 82607 157938 82649 158174
rect 82329 157854 82649 157938
rect 82329 157618 82371 157854
rect 82607 157618 82649 157854
rect 82329 157586 82649 157618
rect 90171 158174 90491 158206
rect 90171 157938 90213 158174
rect 90449 157938 90491 158174
rect 90171 157854 90491 157938
rect 90171 157618 90213 157854
rect 90449 157618 90491 157854
rect 90171 157586 90491 157618
rect 98013 158174 98333 158206
rect 98013 157938 98055 158174
rect 98291 157938 98333 158174
rect 98013 157854 98333 157938
rect 98013 157618 98055 157854
rect 98291 157618 98333 157854
rect 98013 157586 98333 157618
rect 105855 158174 106175 158206
rect 105855 157938 105897 158174
rect 106133 157938 106175 158174
rect 105855 157854 106175 157938
rect 105855 157618 105897 157854
rect 106133 157618 106175 157854
rect 105855 157586 106175 157618
rect 149936 158174 150256 158206
rect 149936 157938 149978 158174
rect 150214 157938 150256 158174
rect 149936 157854 150256 157938
rect 149936 157618 149978 157854
rect 150214 157618 150256 157854
rect 149936 157586 150256 157618
rect 180656 158174 180976 158206
rect 180656 157938 180698 158174
rect 180934 157938 180976 158174
rect 180656 157854 180976 157938
rect 180656 157618 180698 157854
rect 180934 157618 180976 157854
rect 180656 157586 180976 157618
rect 277220 158174 277540 158206
rect 277220 157938 277262 158174
rect 277498 157938 277540 158174
rect 277220 157854 277540 157938
rect 277220 157618 277262 157854
rect 277498 157618 277540 157854
rect 277220 157586 277540 157618
rect 52118 154454 52438 154486
rect 52118 154218 52160 154454
rect 52396 154218 52438 154454
rect 52118 154134 52438 154218
rect 52118 153898 52160 154134
rect 52396 153898 52438 154134
rect 52118 153866 52438 153898
rect 59960 154454 60280 154486
rect 59960 154218 60002 154454
rect 60238 154218 60280 154454
rect 59960 154134 60280 154218
rect 59960 153898 60002 154134
rect 60238 153898 60280 154134
rect 59960 153866 60280 153898
rect 67802 154454 68122 154486
rect 67802 154218 67844 154454
rect 68080 154218 68122 154454
rect 67802 154134 68122 154218
rect 67802 153898 67844 154134
rect 68080 153898 68122 154134
rect 67802 153866 68122 153898
rect 75644 154454 75964 154486
rect 75644 154218 75686 154454
rect 75922 154218 75964 154454
rect 75644 154134 75964 154218
rect 75644 153898 75686 154134
rect 75922 153898 75964 154134
rect 75644 153866 75964 153898
rect 86250 154454 86570 154486
rect 86250 154218 86292 154454
rect 86528 154218 86570 154454
rect 86250 154134 86570 154218
rect 86250 153898 86292 154134
rect 86528 153898 86570 154134
rect 86250 153866 86570 153898
rect 94092 154454 94412 154486
rect 94092 154218 94134 154454
rect 94370 154218 94412 154454
rect 94092 154134 94412 154218
rect 94092 153898 94134 154134
rect 94370 153898 94412 154134
rect 94092 153866 94412 153898
rect 101934 154454 102254 154486
rect 101934 154218 101976 154454
rect 102212 154218 102254 154454
rect 101934 154134 102254 154218
rect 101934 153898 101976 154134
rect 102212 153898 102254 154134
rect 101934 153866 102254 153898
rect 109776 154454 110096 154486
rect 109776 154218 109818 154454
rect 110054 154218 110096 154454
rect 109776 154134 110096 154218
rect 109776 153898 109818 154134
rect 110054 153898 110096 154134
rect 109776 153866 110096 153898
rect 165296 154454 165616 154486
rect 165296 154218 165338 154454
rect 165574 154218 165616 154454
rect 165296 154134 165616 154218
rect 165296 153898 165338 154134
rect 165574 153898 165616 154134
rect 165296 153866 165616 153898
rect 277772 154454 278092 154486
rect 277772 154218 277814 154454
rect 278050 154218 278092 154454
rect 277772 154134 278092 154218
rect 277772 153898 277814 154134
rect 278050 153898 278092 154134
rect 277772 153866 278092 153898
rect 48197 148174 48517 148206
rect 48197 147938 48239 148174
rect 48475 147938 48517 148174
rect 48197 147854 48517 147938
rect 48197 147618 48239 147854
rect 48475 147618 48517 147854
rect 48197 147586 48517 147618
rect 56039 148174 56359 148206
rect 56039 147938 56081 148174
rect 56317 147938 56359 148174
rect 56039 147854 56359 147938
rect 56039 147618 56081 147854
rect 56317 147618 56359 147854
rect 56039 147586 56359 147618
rect 63881 148174 64201 148206
rect 63881 147938 63923 148174
rect 64159 147938 64201 148174
rect 63881 147854 64201 147938
rect 63881 147618 63923 147854
rect 64159 147618 64201 147854
rect 63881 147586 64201 147618
rect 71723 148174 72043 148206
rect 71723 147938 71765 148174
rect 72001 147938 72043 148174
rect 71723 147854 72043 147938
rect 71723 147618 71765 147854
rect 72001 147618 72043 147854
rect 71723 147586 72043 147618
rect 82329 148174 82649 148206
rect 82329 147938 82371 148174
rect 82607 147938 82649 148174
rect 82329 147854 82649 147938
rect 82329 147618 82371 147854
rect 82607 147618 82649 147854
rect 82329 147586 82649 147618
rect 90171 148174 90491 148206
rect 90171 147938 90213 148174
rect 90449 147938 90491 148174
rect 90171 147854 90491 147938
rect 90171 147618 90213 147854
rect 90449 147618 90491 147854
rect 90171 147586 90491 147618
rect 98013 148174 98333 148206
rect 98013 147938 98055 148174
rect 98291 147938 98333 148174
rect 98013 147854 98333 147938
rect 98013 147618 98055 147854
rect 98291 147618 98333 147854
rect 98013 147586 98333 147618
rect 105855 148174 106175 148206
rect 105855 147938 105897 148174
rect 106133 147938 106175 148174
rect 105855 147854 106175 147938
rect 105855 147618 105897 147854
rect 106133 147618 106175 147854
rect 105855 147586 106175 147618
rect 149936 148174 150256 148206
rect 149936 147938 149978 148174
rect 150214 147938 150256 148174
rect 149936 147854 150256 147938
rect 149936 147618 149978 147854
rect 150214 147618 150256 147854
rect 149936 147586 150256 147618
rect 180656 148174 180976 148206
rect 180656 147938 180698 148174
rect 180934 147938 180976 148174
rect 180656 147854 180976 147938
rect 180656 147618 180698 147854
rect 180934 147618 180976 147854
rect 180656 147586 180976 147618
rect 277220 148174 277540 148206
rect 277220 147938 277262 148174
rect 277498 147938 277540 148174
rect 277220 147854 277540 147938
rect 277220 147618 277262 147854
rect 277498 147618 277540 147854
rect 277220 147586 277540 147618
rect 52118 144454 52438 144486
rect 52118 144218 52160 144454
rect 52396 144218 52438 144454
rect 52118 144134 52438 144218
rect 52118 143898 52160 144134
rect 52396 143898 52438 144134
rect 52118 143866 52438 143898
rect 59960 144454 60280 144486
rect 59960 144218 60002 144454
rect 60238 144218 60280 144454
rect 59960 144134 60280 144218
rect 59960 143898 60002 144134
rect 60238 143898 60280 144134
rect 59960 143866 60280 143898
rect 67802 144454 68122 144486
rect 67802 144218 67844 144454
rect 68080 144218 68122 144454
rect 67802 144134 68122 144218
rect 67802 143898 67844 144134
rect 68080 143898 68122 144134
rect 67802 143866 68122 143898
rect 75644 144454 75964 144486
rect 75644 144218 75686 144454
rect 75922 144218 75964 144454
rect 75644 144134 75964 144218
rect 75644 143898 75686 144134
rect 75922 143898 75964 144134
rect 75644 143866 75964 143898
rect 86250 144454 86570 144486
rect 86250 144218 86292 144454
rect 86528 144218 86570 144454
rect 86250 144134 86570 144218
rect 86250 143898 86292 144134
rect 86528 143898 86570 144134
rect 86250 143866 86570 143898
rect 94092 144454 94412 144486
rect 94092 144218 94134 144454
rect 94370 144218 94412 144454
rect 94092 144134 94412 144218
rect 94092 143898 94134 144134
rect 94370 143898 94412 144134
rect 94092 143866 94412 143898
rect 101934 144454 102254 144486
rect 101934 144218 101976 144454
rect 102212 144218 102254 144454
rect 101934 144134 102254 144218
rect 101934 143898 101976 144134
rect 102212 143898 102254 144134
rect 101934 143866 102254 143898
rect 109776 144454 110096 144486
rect 109776 144218 109818 144454
rect 110054 144218 110096 144454
rect 109776 144134 110096 144218
rect 109776 143898 109818 144134
rect 110054 143898 110096 144134
rect 109776 143866 110096 143898
rect 165296 144454 165616 144486
rect 165296 144218 165338 144454
rect 165574 144218 165616 144454
rect 165296 144134 165616 144218
rect 165296 143898 165338 144134
rect 165574 143898 165616 144134
rect 165296 143866 165616 143898
rect 277772 144454 278092 144486
rect 277772 144218 277814 144454
rect 278050 144218 278092 144454
rect 277772 144134 278092 144218
rect 277772 143898 277814 144134
rect 278050 143898 278092 144134
rect 277772 143866 278092 143898
rect 48197 138174 48517 138206
rect 48197 137938 48239 138174
rect 48475 137938 48517 138174
rect 48197 137854 48517 137938
rect 48197 137618 48239 137854
rect 48475 137618 48517 137854
rect 48197 137586 48517 137618
rect 56039 138174 56359 138206
rect 56039 137938 56081 138174
rect 56317 137938 56359 138174
rect 56039 137854 56359 137938
rect 56039 137618 56081 137854
rect 56317 137618 56359 137854
rect 56039 137586 56359 137618
rect 63881 138174 64201 138206
rect 63881 137938 63923 138174
rect 64159 137938 64201 138174
rect 63881 137854 64201 137938
rect 63881 137618 63923 137854
rect 64159 137618 64201 137854
rect 63881 137586 64201 137618
rect 71723 138174 72043 138206
rect 71723 137938 71765 138174
rect 72001 137938 72043 138174
rect 71723 137854 72043 137938
rect 71723 137618 71765 137854
rect 72001 137618 72043 137854
rect 71723 137586 72043 137618
rect 82329 138174 82649 138206
rect 82329 137938 82371 138174
rect 82607 137938 82649 138174
rect 82329 137854 82649 137938
rect 82329 137618 82371 137854
rect 82607 137618 82649 137854
rect 82329 137586 82649 137618
rect 90171 138174 90491 138206
rect 90171 137938 90213 138174
rect 90449 137938 90491 138174
rect 90171 137854 90491 137938
rect 90171 137618 90213 137854
rect 90449 137618 90491 137854
rect 90171 137586 90491 137618
rect 98013 138174 98333 138206
rect 98013 137938 98055 138174
rect 98291 137938 98333 138174
rect 98013 137854 98333 137938
rect 98013 137618 98055 137854
rect 98291 137618 98333 137854
rect 98013 137586 98333 137618
rect 105855 138174 106175 138206
rect 105855 137938 105897 138174
rect 106133 137938 106175 138174
rect 105855 137854 106175 137938
rect 105855 137618 105897 137854
rect 106133 137618 106175 137854
rect 105855 137586 106175 137618
rect 149936 138174 150256 138206
rect 149936 137938 149978 138174
rect 150214 137938 150256 138174
rect 149936 137854 150256 137938
rect 149936 137618 149978 137854
rect 150214 137618 150256 137854
rect 149936 137586 150256 137618
rect 180656 138174 180976 138206
rect 180656 137938 180698 138174
rect 180934 137938 180976 138174
rect 180656 137854 180976 137938
rect 180656 137618 180698 137854
rect 180934 137618 180976 137854
rect 180656 137586 180976 137618
rect 211376 138174 211696 138206
rect 211376 137938 211418 138174
rect 211654 137938 211696 138174
rect 211376 137854 211696 137938
rect 211376 137618 211418 137854
rect 211654 137618 211696 137854
rect 211376 137586 211696 137618
rect 242096 138174 242416 138206
rect 242096 137938 242138 138174
rect 242374 137938 242416 138174
rect 242096 137854 242416 137938
rect 242096 137618 242138 137854
rect 242374 137618 242416 137854
rect 242096 137586 242416 137618
rect 272816 138174 273136 138206
rect 272816 137938 272858 138174
rect 273094 137938 273136 138174
rect 272816 137854 273136 137938
rect 272816 137618 272858 137854
rect 273094 137618 273136 137854
rect 272816 137586 273136 137618
rect 277220 138174 277540 138206
rect 277220 137938 277262 138174
rect 277498 137938 277540 138174
rect 277220 137854 277540 137938
rect 277220 137618 277262 137854
rect 277498 137618 277540 137854
rect 277220 137586 277540 137618
rect 13408 128174 13728 128206
rect 13408 127938 13450 128174
rect 13686 127938 13728 128174
rect 13408 127854 13728 127938
rect 13408 127618 13450 127854
rect 13686 127618 13728 127854
rect 13408 127586 13728 127618
rect 44128 128174 44448 128206
rect 44128 127938 44170 128174
rect 44406 127938 44448 128174
rect 44128 127854 44448 127938
rect 44128 127618 44170 127854
rect 44406 127618 44448 127854
rect 44128 127586 44448 127618
rect 74848 128174 75168 128206
rect 74848 127938 74890 128174
rect 75126 127938 75168 128174
rect 74848 127854 75168 127938
rect 74848 127618 74890 127854
rect 75126 127618 75168 127854
rect 74848 127586 75168 127618
rect 105568 128174 105888 128206
rect 105568 127938 105610 128174
rect 105846 127938 105888 128174
rect 105568 127854 105888 127938
rect 105568 127618 105610 127854
rect 105846 127618 105888 127854
rect 105568 127586 105888 127618
rect 136288 128174 136608 128206
rect 136288 127938 136330 128174
rect 136566 127938 136608 128174
rect 136288 127854 136608 127938
rect 136288 127618 136330 127854
rect 136566 127618 136608 127854
rect 136288 127586 136608 127618
rect 167008 128174 167328 128206
rect 167008 127938 167050 128174
rect 167286 127938 167328 128174
rect 167008 127854 167328 127938
rect 167008 127618 167050 127854
rect 167286 127618 167328 127854
rect 167008 127586 167328 127618
rect 197728 128174 198048 128206
rect 197728 127938 197770 128174
rect 198006 127938 198048 128174
rect 197728 127854 198048 127938
rect 197728 127618 197770 127854
rect 198006 127618 198048 127854
rect 197728 127586 198048 127618
rect 228448 128174 228768 128206
rect 228448 127938 228490 128174
rect 228726 127938 228768 128174
rect 228448 127854 228768 127938
rect 228448 127618 228490 127854
rect 228726 127618 228768 127854
rect 228448 127586 228768 127618
rect 259168 128174 259488 128206
rect 259168 127938 259210 128174
rect 259446 127938 259488 128174
rect 259168 127854 259488 127938
rect 259168 127618 259210 127854
rect 259446 127618 259488 127854
rect 259168 127586 259488 127618
rect 28768 124454 29088 124486
rect 28768 124218 28810 124454
rect 29046 124218 29088 124454
rect 28768 124134 29088 124218
rect 28768 123898 28810 124134
rect 29046 123898 29088 124134
rect 28768 123866 29088 123898
rect 59488 124454 59808 124486
rect 59488 124218 59530 124454
rect 59766 124218 59808 124454
rect 59488 124134 59808 124218
rect 59488 123898 59530 124134
rect 59766 123898 59808 124134
rect 59488 123866 59808 123898
rect 90208 124454 90528 124486
rect 90208 124218 90250 124454
rect 90486 124218 90528 124454
rect 90208 124134 90528 124218
rect 90208 123898 90250 124134
rect 90486 123898 90528 124134
rect 90208 123866 90528 123898
rect 120928 124454 121248 124486
rect 120928 124218 120970 124454
rect 121206 124218 121248 124454
rect 120928 124134 121248 124218
rect 120928 123898 120970 124134
rect 121206 123898 121248 124134
rect 120928 123866 121248 123898
rect 151648 124454 151968 124486
rect 151648 124218 151690 124454
rect 151926 124218 151968 124454
rect 151648 124134 151968 124218
rect 151648 123898 151690 124134
rect 151926 123898 151968 124134
rect 151648 123866 151968 123898
rect 182368 124454 182688 124486
rect 182368 124218 182410 124454
rect 182646 124218 182688 124454
rect 182368 124134 182688 124218
rect 182368 123898 182410 124134
rect 182646 123898 182688 124134
rect 182368 123866 182688 123898
rect 213088 124454 213408 124486
rect 213088 124218 213130 124454
rect 213366 124218 213408 124454
rect 213088 124134 213408 124218
rect 213088 123898 213130 124134
rect 213366 123898 213408 124134
rect 213088 123866 213408 123898
rect 243808 124454 244128 124486
rect 243808 124218 243850 124454
rect 244086 124218 244128 124454
rect 243808 124134 244128 124218
rect 243808 123898 243850 124134
rect 244086 123898 244128 124134
rect 243808 123866 244128 123898
rect 274528 124454 274848 124486
rect 274528 124218 274570 124454
rect 274806 124218 274848 124454
rect 274528 124134 274848 124218
rect 274528 123898 274570 124134
rect 274806 123898 274848 124134
rect 274528 123866 274848 123898
rect 13408 118174 13728 118206
rect 13408 117938 13450 118174
rect 13686 117938 13728 118174
rect 13408 117854 13728 117938
rect 13408 117618 13450 117854
rect 13686 117618 13728 117854
rect 13408 117586 13728 117618
rect 44128 118174 44448 118206
rect 44128 117938 44170 118174
rect 44406 117938 44448 118174
rect 44128 117854 44448 117938
rect 44128 117618 44170 117854
rect 44406 117618 44448 117854
rect 44128 117586 44448 117618
rect 74848 118174 75168 118206
rect 74848 117938 74890 118174
rect 75126 117938 75168 118174
rect 74848 117854 75168 117938
rect 74848 117618 74890 117854
rect 75126 117618 75168 117854
rect 74848 117586 75168 117618
rect 105568 118174 105888 118206
rect 105568 117938 105610 118174
rect 105846 117938 105888 118174
rect 105568 117854 105888 117938
rect 105568 117618 105610 117854
rect 105846 117618 105888 117854
rect 105568 117586 105888 117618
rect 136288 118174 136608 118206
rect 136288 117938 136330 118174
rect 136566 117938 136608 118174
rect 136288 117854 136608 117938
rect 136288 117618 136330 117854
rect 136566 117618 136608 117854
rect 136288 117586 136608 117618
rect 167008 118174 167328 118206
rect 167008 117938 167050 118174
rect 167286 117938 167328 118174
rect 167008 117854 167328 117938
rect 167008 117618 167050 117854
rect 167286 117618 167328 117854
rect 167008 117586 167328 117618
rect 197728 118174 198048 118206
rect 197728 117938 197770 118174
rect 198006 117938 198048 118174
rect 197728 117854 198048 117938
rect 197728 117618 197770 117854
rect 198006 117618 198048 117854
rect 197728 117586 198048 117618
rect 228448 118174 228768 118206
rect 228448 117938 228490 118174
rect 228726 117938 228768 118174
rect 228448 117854 228768 117938
rect 228448 117618 228490 117854
rect 228726 117618 228768 117854
rect 228448 117586 228768 117618
rect 259168 118174 259488 118206
rect 259168 117938 259210 118174
rect 259446 117938 259488 118174
rect 259168 117854 259488 117938
rect 259168 117618 259210 117854
rect 259446 117618 259488 117854
rect 259168 117586 259488 117618
rect 28768 114454 29088 114486
rect 28768 114218 28810 114454
rect 29046 114218 29088 114454
rect 28768 114134 29088 114218
rect 28768 113898 28810 114134
rect 29046 113898 29088 114134
rect 28768 113866 29088 113898
rect 59488 114454 59808 114486
rect 59488 114218 59530 114454
rect 59766 114218 59808 114454
rect 59488 114134 59808 114218
rect 59488 113898 59530 114134
rect 59766 113898 59808 114134
rect 59488 113866 59808 113898
rect 90208 114454 90528 114486
rect 90208 114218 90250 114454
rect 90486 114218 90528 114454
rect 90208 114134 90528 114218
rect 90208 113898 90250 114134
rect 90486 113898 90528 114134
rect 90208 113866 90528 113898
rect 120928 114454 121248 114486
rect 120928 114218 120970 114454
rect 121206 114218 121248 114454
rect 120928 114134 121248 114218
rect 120928 113898 120970 114134
rect 121206 113898 121248 114134
rect 120928 113866 121248 113898
rect 151648 114454 151968 114486
rect 151648 114218 151690 114454
rect 151926 114218 151968 114454
rect 151648 114134 151968 114218
rect 151648 113898 151690 114134
rect 151926 113898 151968 114134
rect 151648 113866 151968 113898
rect 182368 114454 182688 114486
rect 182368 114218 182410 114454
rect 182646 114218 182688 114454
rect 182368 114134 182688 114218
rect 182368 113898 182410 114134
rect 182646 113898 182688 114134
rect 182368 113866 182688 113898
rect 213088 114454 213408 114486
rect 213088 114218 213130 114454
rect 213366 114218 213408 114454
rect 213088 114134 213408 114218
rect 213088 113898 213130 114134
rect 213366 113898 213408 114134
rect 213088 113866 213408 113898
rect 243808 114454 244128 114486
rect 243808 114218 243850 114454
rect 244086 114218 244128 114454
rect 243808 114134 244128 114218
rect 243808 113898 243850 114134
rect 244086 113898 244128 114134
rect 243808 113866 244128 113898
rect 274528 114454 274848 114486
rect 274528 114218 274570 114454
rect 274806 114218 274848 114454
rect 274528 114134 274848 114218
rect 274528 113898 274570 114134
rect 274806 113898 274848 114134
rect 274528 113866 274848 113898
rect 13408 108174 13728 108206
rect 13408 107938 13450 108174
rect 13686 107938 13728 108174
rect 13408 107854 13728 107938
rect 13408 107618 13450 107854
rect 13686 107618 13728 107854
rect 13408 107586 13728 107618
rect 44128 108174 44448 108206
rect 44128 107938 44170 108174
rect 44406 107938 44448 108174
rect 44128 107854 44448 107938
rect 44128 107618 44170 107854
rect 44406 107618 44448 107854
rect 44128 107586 44448 107618
rect 74848 108174 75168 108206
rect 74848 107938 74890 108174
rect 75126 107938 75168 108174
rect 74848 107854 75168 107938
rect 74848 107618 74890 107854
rect 75126 107618 75168 107854
rect 74848 107586 75168 107618
rect 105568 108174 105888 108206
rect 105568 107938 105610 108174
rect 105846 107938 105888 108174
rect 105568 107854 105888 107938
rect 105568 107618 105610 107854
rect 105846 107618 105888 107854
rect 105568 107586 105888 107618
rect 136288 108174 136608 108206
rect 136288 107938 136330 108174
rect 136566 107938 136608 108174
rect 136288 107854 136608 107938
rect 136288 107618 136330 107854
rect 136566 107618 136608 107854
rect 136288 107586 136608 107618
rect 167008 108174 167328 108206
rect 167008 107938 167050 108174
rect 167286 107938 167328 108174
rect 167008 107854 167328 107938
rect 167008 107618 167050 107854
rect 167286 107618 167328 107854
rect 167008 107586 167328 107618
rect 197728 108174 198048 108206
rect 197728 107938 197770 108174
rect 198006 107938 198048 108174
rect 197728 107854 198048 107938
rect 197728 107618 197770 107854
rect 198006 107618 198048 107854
rect 197728 107586 198048 107618
rect 228448 108174 228768 108206
rect 228448 107938 228490 108174
rect 228726 107938 228768 108174
rect 228448 107854 228768 107938
rect 228448 107618 228490 107854
rect 228726 107618 228768 107854
rect 228448 107586 228768 107618
rect 259168 108174 259488 108206
rect 259168 107938 259210 108174
rect 259446 107938 259488 108174
rect 259168 107854 259488 107938
rect 259168 107618 259210 107854
rect 259446 107618 259488 107854
rect 259168 107586 259488 107618
rect 28768 104454 29088 104486
rect 28768 104218 28810 104454
rect 29046 104218 29088 104454
rect 28768 104134 29088 104218
rect 28768 103898 28810 104134
rect 29046 103898 29088 104134
rect 28768 103866 29088 103898
rect 59488 104454 59808 104486
rect 59488 104218 59530 104454
rect 59766 104218 59808 104454
rect 59488 104134 59808 104218
rect 59488 103898 59530 104134
rect 59766 103898 59808 104134
rect 59488 103866 59808 103898
rect 90208 104454 90528 104486
rect 90208 104218 90250 104454
rect 90486 104218 90528 104454
rect 90208 104134 90528 104218
rect 90208 103898 90250 104134
rect 90486 103898 90528 104134
rect 90208 103866 90528 103898
rect 120928 104454 121248 104486
rect 120928 104218 120970 104454
rect 121206 104218 121248 104454
rect 120928 104134 121248 104218
rect 120928 103898 120970 104134
rect 121206 103898 121248 104134
rect 120928 103866 121248 103898
rect 151648 104454 151968 104486
rect 151648 104218 151690 104454
rect 151926 104218 151968 104454
rect 151648 104134 151968 104218
rect 151648 103898 151690 104134
rect 151926 103898 151968 104134
rect 151648 103866 151968 103898
rect 182368 104454 182688 104486
rect 182368 104218 182410 104454
rect 182646 104218 182688 104454
rect 182368 104134 182688 104218
rect 182368 103898 182410 104134
rect 182646 103898 182688 104134
rect 182368 103866 182688 103898
rect 213088 104454 213408 104486
rect 213088 104218 213130 104454
rect 213366 104218 213408 104454
rect 213088 104134 213408 104218
rect 213088 103898 213130 104134
rect 213366 103898 213408 104134
rect 213088 103866 213408 103898
rect 243808 104454 244128 104486
rect 243808 104218 243850 104454
rect 244086 104218 244128 104454
rect 243808 104134 244128 104218
rect 243808 103898 243850 104134
rect 244086 103898 244128 104134
rect 243808 103866 244128 103898
rect 274528 104454 274848 104486
rect 274528 104218 274570 104454
rect 274806 104218 274848 104454
rect 274528 104134 274848 104218
rect 274528 103898 274570 104134
rect 274806 103898 274848 104134
rect 274528 103866 274848 103898
rect 13408 98174 13728 98206
rect 13408 97938 13450 98174
rect 13686 97938 13728 98174
rect 13408 97854 13728 97938
rect 13408 97618 13450 97854
rect 13686 97618 13728 97854
rect 13408 97586 13728 97618
rect 44128 98174 44448 98206
rect 44128 97938 44170 98174
rect 44406 97938 44448 98174
rect 44128 97854 44448 97938
rect 44128 97618 44170 97854
rect 44406 97618 44448 97854
rect 44128 97586 44448 97618
rect 74848 98174 75168 98206
rect 74848 97938 74890 98174
rect 75126 97938 75168 98174
rect 74848 97854 75168 97938
rect 74848 97618 74890 97854
rect 75126 97618 75168 97854
rect 74848 97586 75168 97618
rect 105568 98174 105888 98206
rect 105568 97938 105610 98174
rect 105846 97938 105888 98174
rect 105568 97854 105888 97938
rect 105568 97618 105610 97854
rect 105846 97618 105888 97854
rect 105568 97586 105888 97618
rect 136288 98174 136608 98206
rect 136288 97938 136330 98174
rect 136566 97938 136608 98174
rect 136288 97854 136608 97938
rect 136288 97618 136330 97854
rect 136566 97618 136608 97854
rect 136288 97586 136608 97618
rect 167008 98174 167328 98206
rect 167008 97938 167050 98174
rect 167286 97938 167328 98174
rect 167008 97854 167328 97938
rect 167008 97618 167050 97854
rect 167286 97618 167328 97854
rect 167008 97586 167328 97618
rect 197728 98174 198048 98206
rect 197728 97938 197770 98174
rect 198006 97938 198048 98174
rect 197728 97854 198048 97938
rect 197728 97618 197770 97854
rect 198006 97618 198048 97854
rect 197728 97586 198048 97618
rect 228448 98174 228768 98206
rect 228448 97938 228490 98174
rect 228726 97938 228768 98174
rect 228448 97854 228768 97938
rect 228448 97618 228490 97854
rect 228726 97618 228768 97854
rect 228448 97586 228768 97618
rect 259168 98174 259488 98206
rect 259168 97938 259210 98174
rect 259446 97938 259488 98174
rect 259168 97854 259488 97938
rect 259168 97618 259210 97854
rect 259446 97618 259488 97854
rect 259168 97586 259488 97618
rect 28768 94454 29088 94486
rect 28768 94218 28810 94454
rect 29046 94218 29088 94454
rect 28768 94134 29088 94218
rect 28768 93898 28810 94134
rect 29046 93898 29088 94134
rect 28768 93866 29088 93898
rect 59488 94454 59808 94486
rect 59488 94218 59530 94454
rect 59766 94218 59808 94454
rect 59488 94134 59808 94218
rect 59488 93898 59530 94134
rect 59766 93898 59808 94134
rect 59488 93866 59808 93898
rect 90208 94454 90528 94486
rect 90208 94218 90250 94454
rect 90486 94218 90528 94454
rect 90208 94134 90528 94218
rect 90208 93898 90250 94134
rect 90486 93898 90528 94134
rect 90208 93866 90528 93898
rect 120928 94454 121248 94486
rect 120928 94218 120970 94454
rect 121206 94218 121248 94454
rect 120928 94134 121248 94218
rect 120928 93898 120970 94134
rect 121206 93898 121248 94134
rect 120928 93866 121248 93898
rect 151648 94454 151968 94486
rect 151648 94218 151690 94454
rect 151926 94218 151968 94454
rect 151648 94134 151968 94218
rect 151648 93898 151690 94134
rect 151926 93898 151968 94134
rect 151648 93866 151968 93898
rect 182368 94454 182688 94486
rect 182368 94218 182410 94454
rect 182646 94218 182688 94454
rect 182368 94134 182688 94218
rect 182368 93898 182410 94134
rect 182646 93898 182688 94134
rect 182368 93866 182688 93898
rect 213088 94454 213408 94486
rect 213088 94218 213130 94454
rect 213366 94218 213408 94454
rect 213088 94134 213408 94218
rect 213088 93898 213130 94134
rect 213366 93898 213408 94134
rect 213088 93866 213408 93898
rect 243808 94454 244128 94486
rect 243808 94218 243850 94454
rect 244086 94218 244128 94454
rect 243808 94134 244128 94218
rect 243808 93898 243850 94134
rect 244086 93898 244128 94134
rect 243808 93866 244128 93898
rect 274528 94454 274848 94486
rect 274528 94218 274570 94454
rect 274806 94218 274848 94454
rect 274528 94134 274848 94218
rect 274528 93898 274570 94134
rect 274806 93898 274848 94134
rect 274528 93866 274848 93898
rect 274219 89044 274285 89045
rect 274219 88980 274220 89044
rect 274284 88980 274285 89044
rect 274219 88979 274285 88980
rect 272379 87548 272445 87549
rect 272379 87484 272380 87548
rect 272444 87484 272445 87548
rect 272379 87483 272445 87484
rect 9443 21860 9509 21861
rect 9443 21796 9444 21860
rect 9508 21796 9509 21860
rect 9443 21795 9509 21796
rect 272382 19141 272442 87483
rect 273851 76532 273917 76533
rect 273851 76468 273852 76532
rect 273916 76468 273917 76532
rect 273851 76467 273917 76468
rect 272563 65516 272629 65517
rect 272563 65452 272564 65516
rect 272628 65452 272629 65516
rect 272563 65451 272629 65452
rect 272566 20637 272626 65451
rect 273299 22676 273365 22677
rect 273299 22612 273300 22676
rect 273364 22612 273365 22676
rect 273299 22611 273365 22612
rect 272563 20636 272629 20637
rect 272563 20572 272564 20636
rect 272628 20572 272629 20636
rect 272563 20571 272629 20572
rect 273302 20229 273362 22611
rect 273299 20228 273365 20229
rect 273299 20164 273300 20228
rect 273364 20164 273365 20228
rect 273299 20163 273365 20164
rect 273854 19277 273914 76467
rect 274035 66468 274101 66469
rect 274035 66404 274036 66468
rect 274100 66404 274101 66468
rect 274035 66403 274101 66404
rect 274038 62797 274098 66403
rect 274222 65620 274282 88979
rect 278267 86188 278333 86189
rect 278267 86124 278268 86188
rect 278332 86124 278333 86188
rect 278267 86123 278333 86124
rect 277163 84828 277229 84829
rect 277163 84764 277164 84828
rect 277228 84764 277229 84828
rect 277163 84763 277229 84764
rect 276059 83468 276125 83469
rect 276059 83404 276060 83468
rect 276124 83404 276125 83468
rect 276059 83403 276125 83404
rect 274955 77892 275021 77893
rect 274955 77828 274956 77892
rect 275020 77828 275021 77892
rect 274955 77827 275021 77828
rect 274587 68236 274653 68237
rect 274587 68172 274588 68236
rect 274652 68172 274653 68236
rect 274587 68171 274653 68172
rect 274590 65620 274650 68171
rect 274958 65620 275018 77827
rect 275323 75172 275389 75173
rect 275323 75108 275324 75172
rect 275388 75108 275389 75172
rect 275323 75107 275389 75108
rect 275326 65620 275386 75107
rect 275691 68372 275757 68373
rect 275691 68308 275692 68372
rect 275756 68308 275757 68372
rect 275691 68307 275757 68308
rect 275694 65620 275754 68307
rect 276062 65620 276122 83403
rect 276795 82108 276861 82109
rect 276795 82044 276796 82108
rect 276860 82044 276861 82108
rect 276795 82043 276861 82044
rect 276427 73812 276493 73813
rect 276427 73748 276428 73812
rect 276492 73748 276493 73812
rect 276427 73747 276493 73748
rect 276430 65620 276490 73747
rect 276798 65620 276858 82043
rect 277166 65620 277226 84763
rect 277899 80748 277965 80749
rect 277899 80684 277900 80748
rect 277964 80684 277965 80748
rect 277899 80683 277965 80684
rect 277531 72452 277597 72453
rect 277531 72388 277532 72452
rect 277596 72388 277597 72452
rect 277531 72387 277597 72388
rect 277534 65620 277594 72387
rect 277902 65620 277962 80683
rect 278270 65620 278330 86123
rect 278635 67012 278701 67013
rect 278635 66948 278636 67012
rect 278700 66948 278701 67012
rect 278635 66947 278701 66948
rect 278638 65620 278698 66947
rect 279006 65620 279066 179147
rect 281030 178941 281090 182411
rect 281579 181660 281645 181661
rect 281579 181596 281580 181660
rect 281644 181596 281645 181660
rect 281579 181595 281645 181596
rect 281582 181386 281642 181595
rect 281214 181326 281642 181386
rect 281027 178940 281093 178941
rect 281027 178876 281028 178940
rect 281092 178876 281093 178940
rect 281027 178875 281093 178876
rect 280291 178260 280357 178261
rect 280291 178196 280292 178260
rect 280356 178196 280357 178260
rect 280291 178195 280357 178196
rect 279555 175404 279621 175405
rect 279555 175340 279556 175404
rect 279620 175340 279621 175404
rect 279555 175339 279621 175340
rect 279558 68237 279618 175339
rect 280294 74550 280354 178195
rect 281214 177170 281274 181326
rect 281395 180980 281461 180981
rect 281395 180916 281396 180980
rect 281460 180916 281461 180980
rect 281395 180915 281461 180916
rect 281398 177309 281458 180915
rect 281579 180708 281645 180709
rect 281579 180644 281580 180708
rect 281644 180644 281645 180708
rect 281579 180643 281645 180644
rect 281395 177308 281461 177309
rect 281395 177244 281396 177308
rect 281460 177244 281461 177308
rect 281395 177243 281461 177244
rect 281214 177110 281458 177170
rect 281211 176628 281277 176629
rect 281211 176564 281212 176628
rect 281276 176564 281277 176628
rect 281211 176563 281277 176564
rect 280110 74490 280354 74550
rect 279739 69596 279805 69597
rect 279739 69532 279740 69596
rect 279804 69532 279805 69596
rect 279739 69531 279805 69532
rect 279555 68236 279621 68237
rect 279555 68172 279556 68236
rect 279620 68172 279621 68236
rect 279555 68171 279621 68172
rect 279371 66876 279437 66877
rect 279371 66812 279372 66876
rect 279436 66812 279437 66876
rect 279371 66811 279437 66812
rect 279374 65620 279434 66811
rect 279742 65620 279802 69531
rect 280110 65620 280170 74490
rect 281214 65724 281274 176563
rect 281398 157997 281458 177110
rect 281395 157996 281461 157997
rect 281395 157932 281396 157996
rect 281460 157932 281461 157996
rect 281395 157931 281461 157932
rect 281582 65620 281642 180643
rect 281766 179077 281826 214507
rect 281763 179076 281829 179077
rect 281763 179012 281764 179076
rect 281828 179012 281829 179076
rect 281763 179011 281829 179012
rect 281950 175405 282010 281011
rect 284339 280804 284405 280805
rect 284339 280740 284340 280804
rect 284404 280740 284405 280804
rect 284339 280739 284405 280740
rect 282867 190500 282933 190501
rect 282867 190436 282868 190500
rect 282932 190436 282933 190500
rect 282867 190435 282933 190436
rect 282870 190208 282930 190435
rect 282686 190148 282930 190208
rect 282499 189276 282565 189277
rect 282499 189212 282500 189276
rect 282564 189212 282565 189276
rect 282499 189211 282565 189212
rect 282502 184789 282562 189211
rect 282686 186690 282746 190148
rect 283787 189684 283853 189685
rect 283787 189620 283788 189684
rect 283852 189620 283853 189684
rect 283787 189619 283853 189620
rect 283051 189548 283117 189549
rect 283051 189484 283052 189548
rect 283116 189484 283117 189548
rect 283051 189483 283117 189484
rect 282686 186630 282930 186690
rect 282870 186330 282930 186630
rect 282686 186270 282930 186330
rect 282499 184788 282565 184789
rect 282499 184724 282500 184788
rect 282564 184724 282565 184788
rect 282499 184723 282565 184724
rect 282131 184652 282197 184653
rect 282131 184588 282132 184652
rect 282196 184588 282197 184652
rect 282131 184587 282197 184588
rect 282134 180437 282194 184587
rect 282686 184381 282746 186270
rect 282683 184380 282749 184381
rect 282683 184316 282684 184380
rect 282748 184316 282749 184380
rect 282683 184315 282749 184316
rect 283054 181389 283114 189483
rect 283419 187916 283485 187917
rect 283419 187852 283420 187916
rect 283484 187852 283485 187916
rect 283419 187851 283485 187852
rect 283422 184925 283482 187851
rect 283790 187237 283850 189619
rect 283971 189140 284037 189141
rect 283971 189076 283972 189140
rect 284036 189076 284037 189140
rect 283971 189075 284037 189076
rect 283787 187236 283853 187237
rect 283787 187172 283788 187236
rect 283852 187172 283853 187236
rect 283787 187171 283853 187172
rect 283603 186692 283669 186693
rect 283603 186628 283604 186692
rect 283668 186628 283669 186692
rect 283603 186627 283669 186628
rect 283606 186285 283666 186627
rect 283603 186284 283669 186285
rect 283603 186220 283604 186284
rect 283668 186220 283669 186284
rect 283603 186219 283669 186220
rect 283974 186149 284034 189075
rect 284155 188596 284221 188597
rect 284155 188532 284156 188596
rect 284220 188532 284221 188596
rect 284155 188531 284221 188532
rect 283971 186148 284037 186149
rect 283971 186084 283972 186148
rect 284036 186084 284037 186148
rect 283971 186083 284037 186084
rect 284158 186013 284218 188531
rect 284342 186829 284402 280739
rect 284523 193220 284589 193221
rect 284523 193156 284524 193220
rect 284588 193156 284589 193220
rect 284523 193155 284589 193156
rect 284339 186828 284405 186829
rect 284339 186764 284340 186828
rect 284404 186764 284405 186828
rect 284339 186763 284405 186764
rect 284155 186012 284221 186013
rect 284155 185948 284156 186012
rect 284220 185948 284221 186012
rect 284155 185947 284221 185948
rect 283419 184924 283485 184925
rect 283419 184860 283420 184924
rect 283484 184860 283485 184924
rect 283419 184859 283485 184860
rect 284155 181524 284221 181525
rect 284155 181460 284156 181524
rect 284220 181460 284221 181524
rect 284155 181459 284221 181460
rect 283051 181388 283117 181389
rect 283051 181324 283052 181388
rect 283116 181324 283117 181388
rect 283051 181323 283117 181324
rect 283051 181252 283117 181253
rect 283051 181188 283052 181252
rect 283116 181188 283117 181252
rect 283051 181187 283117 181188
rect 282683 180844 282749 180845
rect 282683 180780 282684 180844
rect 282748 180780 282749 180844
rect 282683 180779 282749 180780
rect 282131 180436 282197 180437
rect 282131 180372 282132 180436
rect 282196 180372 282197 180436
rect 282131 180371 282197 180372
rect 282131 177308 282197 177309
rect 282131 177244 282132 177308
rect 282196 177244 282197 177308
rect 282131 177243 282197 177244
rect 281947 175404 282013 175405
rect 281947 175340 281948 175404
rect 282012 175340 282013 175404
rect 281947 175339 282013 175340
rect 281947 175268 282013 175269
rect 281947 175204 281948 175268
rect 282012 175204 282013 175268
rect 281947 175203 282013 175204
rect 281950 65620 282010 175203
rect 282134 171150 282194 177243
rect 282686 177170 282746 180779
rect 282686 177110 282930 177170
rect 282683 176764 282749 176765
rect 282683 176700 282684 176764
rect 282748 176700 282749 176764
rect 282683 176699 282749 176700
rect 282134 171090 282378 171150
rect 282318 65620 282378 171090
rect 282686 65620 282746 176699
rect 282870 175269 282930 177110
rect 282867 175268 282933 175269
rect 282867 175204 282868 175268
rect 282932 175204 282933 175268
rect 282867 175203 282933 175204
rect 283054 65620 283114 181187
rect 284158 156637 284218 181459
rect 284526 179213 284586 193155
rect 285259 182068 285325 182069
rect 285259 182004 285260 182068
rect 285324 182004 285325 182068
rect 285259 182003 285325 182004
rect 284707 181116 284773 181117
rect 284707 181052 284708 181116
rect 284772 181052 284773 181116
rect 284707 181051 284773 181052
rect 284523 179212 284589 179213
rect 284523 179148 284524 179212
rect 284588 179148 284589 179212
rect 284523 179147 284589 179148
rect 284710 176765 284770 181051
rect 284891 178940 284957 178941
rect 284891 178876 284892 178940
rect 284956 178876 284957 178940
rect 284891 178875 284957 178876
rect 284707 176764 284773 176765
rect 284707 176700 284708 176764
rect 284772 176700 284773 176764
rect 284707 176699 284773 176700
rect 284894 157453 284954 178875
rect 284891 157452 284957 157453
rect 284891 157388 284892 157452
rect 284956 157388 284957 157452
rect 284891 157387 284957 157388
rect 284155 156636 284221 156637
rect 284155 156572 284156 156636
rect 284220 156572 284221 156636
rect 284155 156571 284221 156572
rect 284891 155276 284957 155277
rect 284891 155212 284892 155276
rect 284956 155212 284957 155276
rect 284891 155211 284957 155212
rect 283787 71228 283853 71229
rect 283787 71164 283788 71228
rect 283852 71164 283853 71228
rect 283787 71163 283853 71164
rect 283419 68780 283485 68781
rect 283419 68716 283420 68780
rect 283484 68716 283485 68780
rect 283419 68715 283485 68716
rect 283422 65620 283482 68715
rect 283790 65620 283850 71163
rect 284707 69732 284773 69733
rect 284707 69668 284708 69732
rect 284772 69668 284773 69732
rect 284707 69667 284773 69668
rect 284155 69596 284221 69597
rect 284155 69532 284156 69596
rect 284220 69532 284221 69596
rect 284155 69531 284221 69532
rect 284158 65620 284218 69531
rect 284710 65650 284770 69667
rect 284556 65590 284770 65650
rect 284894 65620 284954 155211
rect 285262 65620 285322 182003
rect 285443 181796 285509 181797
rect 285443 181732 285444 181796
rect 285508 181732 285509 181796
rect 285443 181731 285509 181732
rect 285446 69733 285506 181731
rect 285630 178261 285690 671195
rect 290411 658204 290477 658205
rect 290411 658140 290412 658204
rect 290476 658140 290477 658204
rect 290411 658139 290477 658140
rect 287099 280940 287165 280941
rect 287099 280876 287100 280940
rect 287164 280876 287165 280940
rect 287099 280875 287165 280876
rect 285811 188732 285877 188733
rect 285811 188668 285812 188732
rect 285876 188668 285877 188732
rect 285811 188667 285877 188668
rect 285814 182205 285874 188667
rect 287102 184925 287162 280875
rect 287099 184924 287165 184925
rect 287099 184860 287100 184924
rect 287164 184860 287165 184924
rect 287099 184859 287165 184860
rect 290227 183972 290293 183973
rect 290227 183908 290228 183972
rect 290292 183908 290293 183972
rect 290227 183907 290293 183908
rect 289491 183700 289557 183701
rect 289491 183636 289492 183700
rect 289556 183636 289557 183700
rect 289491 183635 289557 183636
rect 288939 183428 289005 183429
rect 288939 183364 288940 183428
rect 289004 183364 289005 183428
rect 288939 183363 289005 183364
rect 288203 183156 288269 183157
rect 288203 183092 288204 183156
rect 288268 183092 288269 183156
rect 288203 183091 288269 183092
rect 287835 183020 287901 183021
rect 287835 182956 287836 183020
rect 287900 182956 287901 183020
rect 287835 182955 287901 182956
rect 287467 182884 287533 182885
rect 287467 182820 287468 182884
rect 287532 182820 287533 182884
rect 287467 182819 287533 182820
rect 287099 182748 287165 182749
rect 287099 182684 287100 182748
rect 287164 182684 287165 182748
rect 287099 182683 287165 182684
rect 285995 182340 286061 182341
rect 285995 182276 285996 182340
rect 286060 182276 286061 182340
rect 285995 182275 286061 182276
rect 285811 182204 285877 182205
rect 285811 182140 285812 182204
rect 285876 182140 285877 182204
rect 285811 182139 285877 182140
rect 285627 178260 285693 178261
rect 285627 178196 285628 178260
rect 285692 178196 285693 178260
rect 285627 178195 285693 178196
rect 285443 69732 285509 69733
rect 285443 69668 285444 69732
rect 285508 69668 285509 69732
rect 285443 69667 285509 69668
rect 285814 65650 285874 182139
rect 285660 65590 285874 65650
rect 285998 65620 286058 182275
rect 286731 179212 286797 179213
rect 286731 179148 286732 179212
rect 286796 179148 286797 179212
rect 286731 179147 286797 179148
rect 286363 157452 286429 157453
rect 286363 157388 286364 157452
rect 286428 157388 286429 157452
rect 286363 157387 286429 157388
rect 286366 65620 286426 157387
rect 286734 65620 286794 179147
rect 287102 65620 287162 182683
rect 287470 65620 287530 182819
rect 287838 65620 287898 182955
rect 288206 65620 288266 183091
rect 288571 182204 288637 182205
rect 288571 182140 288572 182204
rect 288636 182140 288637 182204
rect 288571 182139 288637 182140
rect 288574 65620 288634 182139
rect 288942 65620 289002 183363
rect 289307 183292 289373 183293
rect 289307 183228 289308 183292
rect 289372 183228 289373 183292
rect 289307 183227 289373 183228
rect 289310 65620 289370 183227
rect 289494 180810 289554 183635
rect 289675 183564 289741 183565
rect 289675 183500 289676 183564
rect 289740 183500 289741 183564
rect 289675 183499 289741 183500
rect 289678 183293 289738 183499
rect 289675 183292 289741 183293
rect 289675 183228 289676 183292
rect 289740 183228 289741 183292
rect 289675 183227 289741 183228
rect 289494 180750 289738 180810
rect 289678 65670 289738 180750
rect 290043 179484 290109 179485
rect 290043 179420 290044 179484
rect 290108 179420 290109 179484
rect 290043 179419 290109 179420
rect 290046 65620 290106 179419
rect 290230 65754 290290 183907
rect 290414 69597 290474 658139
rect 291699 190500 291765 190501
rect 291699 190436 291700 190500
rect 291764 190436 291765 190500
rect 291699 190435 291765 190436
rect 291147 188052 291213 188053
rect 291147 187988 291148 188052
rect 291212 187988 291213 188052
rect 291147 187987 291213 187988
rect 290595 183836 290661 183837
rect 290595 183772 290596 183836
rect 290660 183772 290661 183836
rect 290595 183771 290661 183772
rect 290598 180301 290658 183771
rect 290595 180300 290661 180301
rect 290595 180236 290596 180300
rect 290660 180236 290661 180300
rect 290595 180235 290661 180236
rect 290598 179485 290658 180235
rect 290595 179484 290661 179485
rect 290595 179420 290596 179484
rect 290660 179420 290661 179484
rect 290595 179419 290661 179420
rect 291150 174589 291210 187987
rect 291515 184108 291581 184109
rect 291515 184044 291516 184108
rect 291580 184044 291581 184108
rect 291515 184043 291581 184044
rect 291147 174588 291213 174589
rect 291147 174524 291148 174588
rect 291212 174524 291213 174588
rect 291147 174523 291213 174524
rect 290411 69596 290477 69597
rect 290411 69532 290412 69596
rect 290476 69532 290477 69596
rect 290411 69531 290477 69532
rect 290230 65694 290444 65754
rect 291518 65620 291578 184043
rect 291702 179077 291762 190435
rect 292803 189276 292869 189277
rect 292803 189212 292804 189276
rect 292868 189212 292869 189276
rect 292803 189211 292869 189212
rect 292619 187916 292685 187917
rect 292619 187852 292620 187916
rect 292684 187852 292685 187916
rect 292619 187851 292685 187852
rect 292622 184925 292682 187851
rect 292619 184924 292685 184925
rect 292619 184860 292620 184924
rect 292684 184860 292685 184924
rect 292619 184859 292685 184860
rect 292806 184789 292866 189211
rect 292987 188324 293053 188325
rect 292987 188260 292988 188324
rect 293052 188260 293053 188324
rect 292987 188259 293053 188260
rect 292803 184788 292869 184789
rect 292803 184724 292804 184788
rect 292868 184724 292869 184788
rect 292803 184723 292869 184724
rect 292619 184516 292685 184517
rect 292619 184452 292620 184516
rect 292684 184452 292685 184516
rect 292619 184451 292685 184452
rect 291883 183836 291949 183837
rect 291883 183772 291884 183836
rect 291948 183772 291949 183836
rect 291883 183771 291949 183772
rect 291699 179076 291765 179077
rect 291699 179012 291700 179076
rect 291764 179012 291765 179076
rect 291699 179011 291765 179012
rect 291702 178125 291762 179011
rect 291699 178124 291765 178125
rect 291699 178060 291700 178124
rect 291764 178060 291765 178124
rect 291699 178059 291765 178060
rect 291886 65620 291946 183771
rect 292251 178124 292317 178125
rect 292251 178060 292252 178124
rect 292316 178060 292317 178124
rect 292251 178059 292317 178060
rect 292254 65620 292314 178059
rect 292622 65620 292682 184451
rect 292990 180437 293050 188259
rect 296299 185876 296365 185877
rect 296299 185812 296300 185876
rect 296364 185812 296365 185876
rect 296299 185811 296365 185812
rect 295931 185740 295997 185741
rect 295931 185676 295932 185740
rect 295996 185676 295997 185740
rect 295931 185675 295997 185676
rect 295563 185604 295629 185605
rect 295563 185540 295564 185604
rect 295628 185540 295629 185604
rect 295563 185539 295629 185540
rect 295195 185468 295261 185469
rect 295195 185404 295196 185468
rect 295260 185404 295261 185468
rect 295195 185403 295261 185404
rect 294827 185332 294893 185333
rect 294827 185268 294828 185332
rect 294892 185268 294893 185332
rect 294827 185267 294893 185268
rect 294459 185196 294525 185197
rect 294459 185132 294460 185196
rect 294524 185132 294525 185196
rect 294459 185131 294525 185132
rect 294091 185060 294157 185061
rect 294091 184996 294092 185060
rect 294156 184996 294157 185060
rect 294091 184995 294157 184996
rect 293723 184924 293789 184925
rect 293723 184860 293724 184924
rect 293788 184860 293789 184924
rect 293723 184859 293789 184860
rect 293355 184788 293421 184789
rect 293355 184724 293356 184788
rect 293420 184724 293421 184788
rect 293355 184723 293421 184724
rect 292987 180436 293053 180437
rect 292987 180372 292988 180436
rect 293052 180372 293053 180436
rect 292987 180371 293053 180372
rect 292990 65620 293050 180371
rect 293358 65620 293418 184723
rect 293726 65620 293786 184859
rect 294094 65620 294154 184995
rect 294462 65620 294522 185131
rect 294830 65620 294890 185267
rect 295198 65620 295258 185403
rect 295566 65620 295626 185539
rect 295934 65620 295994 185675
rect 296302 178941 296362 185811
rect 296299 178940 296365 178941
rect 296299 178876 296300 178940
rect 296364 178876 296365 178940
rect 296299 178875 296365 178876
rect 296302 65620 296362 178875
rect 296486 156909 296546 700299
rect 585310 698174 585930 704282
rect 585310 697938 585342 698174
rect 585578 697938 585662 698174
rect 585898 697938 585930 698174
rect 585310 697854 585930 697938
rect 585310 697618 585342 697854
rect 585578 697618 585662 697854
rect 585898 697618 585930 697854
rect 585310 688174 585930 697618
rect 585310 687938 585342 688174
rect 585578 687938 585662 688174
rect 585898 687938 585930 688174
rect 585310 687854 585930 687938
rect 585310 687618 585342 687854
rect 585578 687618 585662 687854
rect 585898 687618 585930 687854
rect 585310 678174 585930 687618
rect 585310 677938 585342 678174
rect 585578 677938 585662 678174
rect 585898 677938 585930 678174
rect 585310 677854 585930 677938
rect 585310 677618 585342 677854
rect 585578 677618 585662 677854
rect 585898 677618 585930 677854
rect 575979 670716 576045 670717
rect 575979 670652 575980 670716
rect 576044 670652 576045 670716
rect 575979 670651 576045 670652
rect 574691 564364 574757 564365
rect 574691 564300 574692 564364
rect 574756 564300 574757 564364
rect 574691 564299 574757 564300
rect 420957 323508 421023 323509
rect 420957 323444 420958 323508
rect 421022 323444 421023 323508
rect 420957 323443 421023 323444
rect 422181 323508 422247 323509
rect 422181 323444 422182 323508
rect 422246 323444 422247 323508
rect 422181 323443 422247 323444
rect 433333 323508 433399 323509
rect 433333 323444 433334 323508
rect 433398 323444 433399 323508
rect 433333 323443 433399 323444
rect 420960 323202 421020 323443
rect 422184 323202 422244 323443
rect 433336 323202 433396 323443
rect 441659 319292 441725 319293
rect 441659 319228 441660 319292
rect 441724 319228 441725 319292
rect 441659 319227 441725 319228
rect 303448 318174 303796 318206
rect 303448 317938 303504 318174
rect 303740 317938 303796 318174
rect 303448 317854 303796 317938
rect 303448 317618 303504 317854
rect 303740 317618 303796 317854
rect 303448 317586 303796 317618
rect 437816 318174 438164 318206
rect 437816 317938 437872 318174
rect 438108 317938 438164 318174
rect 437816 317854 438164 317938
rect 437816 317618 437872 317854
rect 438108 317618 438164 317854
rect 437816 317586 438164 317618
rect 302768 314454 303116 314486
rect 302768 314218 302824 314454
rect 303060 314218 303116 314454
rect 302768 314134 303116 314218
rect 302768 313898 302824 314134
rect 303060 313898 303116 314134
rect 302768 313866 303116 313898
rect 438496 314454 438844 314486
rect 438496 314218 438552 314454
rect 438788 314218 438844 314454
rect 438496 314134 438844 314218
rect 438496 313898 438552 314134
rect 438788 313898 438844 314134
rect 438496 313866 438844 313898
rect 303448 308174 303796 308206
rect 303448 307938 303504 308174
rect 303740 307938 303796 308174
rect 303448 307854 303796 307938
rect 303448 307618 303504 307854
rect 303740 307618 303796 307854
rect 303448 307586 303796 307618
rect 437816 308174 438164 308206
rect 437816 307938 437872 308174
rect 438108 307938 438164 308174
rect 437816 307854 438164 307938
rect 437816 307618 437872 307854
rect 438108 307618 438164 307854
rect 437816 307586 438164 307618
rect 302768 304454 303116 304486
rect 302768 304218 302824 304454
rect 303060 304218 303116 304454
rect 302768 304134 303116 304218
rect 302768 303898 302824 304134
rect 303060 303898 303116 304134
rect 302768 303866 303116 303898
rect 438496 304454 438844 304486
rect 438496 304218 438552 304454
rect 438788 304218 438844 304454
rect 438496 304134 438844 304218
rect 438496 303898 438552 304134
rect 438788 303898 438844 304134
rect 438496 303866 438844 303898
rect 303448 298174 303796 298206
rect 303448 297938 303504 298174
rect 303740 297938 303796 298174
rect 303448 297854 303796 297938
rect 303448 297618 303504 297854
rect 303740 297618 303796 297854
rect 303448 297586 303796 297618
rect 437816 298174 438164 298206
rect 437816 297938 437872 298174
rect 438108 297938 438164 298174
rect 437816 297854 438164 297938
rect 437816 297618 437872 297854
rect 438108 297618 438164 297854
rect 437816 297586 438164 297618
rect 302768 294454 303116 294486
rect 302768 294218 302824 294454
rect 303060 294218 303116 294454
rect 302768 294134 303116 294218
rect 302768 293898 302824 294134
rect 303060 293898 303116 294134
rect 302768 293866 303116 293898
rect 438496 294454 438844 294486
rect 438496 294218 438552 294454
rect 438788 294218 438844 294454
rect 438496 294134 438844 294218
rect 438496 293898 438552 294134
rect 438788 293898 438844 294134
rect 438496 293866 438844 293898
rect 303448 288174 303796 288206
rect 303448 287938 303504 288174
rect 303740 287938 303796 288174
rect 303448 287854 303796 287938
rect 303448 287618 303504 287854
rect 303740 287618 303796 287854
rect 303448 287586 303796 287618
rect 437816 288174 438164 288206
rect 437816 287938 437872 288174
rect 438108 287938 438164 288174
rect 437816 287854 438164 287938
rect 437816 287618 437872 287854
rect 438108 287618 438164 287854
rect 437816 287586 438164 287618
rect 302768 284454 303116 284486
rect 302768 284218 302824 284454
rect 303060 284218 303116 284454
rect 302768 284134 303116 284218
rect 302768 283898 302824 284134
rect 303060 283898 303116 284134
rect 302768 283866 303116 283898
rect 438496 284454 438844 284486
rect 438496 284218 438552 284454
rect 438788 284218 438844 284454
rect 438496 284134 438844 284218
rect 438496 283898 438552 284134
rect 438788 283898 438844 284134
rect 438496 283866 438844 283898
rect 303448 278174 303796 278206
rect 303448 277938 303504 278174
rect 303740 277938 303796 278174
rect 303448 277854 303796 277938
rect 303448 277618 303504 277854
rect 303740 277618 303796 277854
rect 303448 277586 303796 277618
rect 437816 278174 438164 278206
rect 437816 277938 437872 278174
rect 438108 277938 438164 278174
rect 437816 277854 438164 277938
rect 437816 277618 437872 277854
rect 438108 277618 438164 277854
rect 437816 277586 438164 277618
rect 300531 276860 300597 276861
rect 300531 276796 300532 276860
rect 300596 276796 300597 276860
rect 300531 276795 300597 276796
rect 300163 269924 300229 269925
rect 300163 269860 300164 269924
rect 300228 269860 300229 269924
rect 300163 269859 300229 269860
rect 299979 248300 300045 248301
rect 299979 248236 299980 248300
rect 300044 248236 300045 248300
rect 299979 248235 300045 248236
rect 299982 236061 300042 248235
rect 300166 247077 300226 269859
rect 300347 268156 300413 268157
rect 300347 268092 300348 268156
rect 300412 268092 300413 268156
rect 300347 268091 300413 268092
rect 300163 247076 300229 247077
rect 300163 247012 300164 247076
rect 300228 247012 300229 247076
rect 300163 247011 300229 247012
rect 300350 237421 300410 268091
rect 300534 249797 300594 276795
rect 302003 275974 302069 275975
rect 302003 275910 302004 275974
rect 302068 275910 302069 275974
rect 302003 275909 302069 275910
rect 301819 273732 301885 273733
rect 301819 273668 301820 273732
rect 301884 273668 301885 273732
rect 301819 273667 301885 273668
rect 301635 272780 301701 272781
rect 301635 272716 301636 272780
rect 301700 272716 301701 272780
rect 301635 272715 301701 272716
rect 300715 271012 300781 271013
rect 300715 270948 300716 271012
rect 300780 270948 300781 271012
rect 300715 270947 300781 270948
rect 300531 249796 300597 249797
rect 300531 249732 300532 249796
rect 300596 249732 300597 249796
rect 300531 249731 300597 249732
rect 300531 248028 300597 248029
rect 300531 247964 300532 248028
rect 300596 247964 300597 248028
rect 300531 247963 300597 247964
rect 300347 237420 300413 237421
rect 300347 237356 300348 237420
rect 300412 237356 300413 237420
rect 300347 237355 300413 237356
rect 299979 236060 300045 236061
rect 299979 235996 299980 236060
rect 300044 235996 300045 236060
rect 299979 235995 300045 235996
rect 300534 217429 300594 247963
rect 300718 235925 300778 270947
rect 301451 249932 301517 249933
rect 301451 249868 301452 249932
rect 301516 249868 301517 249932
rect 301451 249867 301517 249868
rect 301454 240005 301514 249867
rect 301451 240004 301517 240005
rect 301451 239940 301452 240004
rect 301516 239940 301517 240004
rect 301451 239939 301517 239940
rect 300715 235924 300781 235925
rect 300715 235860 300716 235924
rect 300780 235860 300781 235924
rect 300715 235859 300781 235860
rect 301638 233885 301698 272715
rect 301635 233884 301701 233885
rect 301635 233820 301636 233884
rect 301700 233820 301701 233884
rect 301635 233819 301701 233820
rect 301822 232525 301882 273667
rect 301819 232524 301885 232525
rect 301819 232460 301820 232524
rect 301884 232460 301885 232524
rect 301819 232459 301885 232460
rect 302006 218653 302066 275909
rect 302768 274454 303116 274486
rect 302768 274218 302824 274454
rect 303060 274218 303116 274454
rect 302768 274134 303116 274218
rect 302768 273898 302824 274134
rect 303060 273898 303116 274134
rect 302768 273866 303116 273898
rect 438496 274454 438844 274486
rect 438496 274218 438552 274454
rect 438788 274218 438844 274454
rect 438496 274134 438844 274218
rect 438496 273898 438552 274134
rect 438788 273898 438844 274134
rect 438496 273866 438844 273898
rect 303448 268174 303796 268206
rect 303448 267938 303504 268174
rect 303740 267938 303796 268174
rect 303448 267854 303796 267938
rect 303448 267618 303504 267854
rect 303740 267618 303796 267854
rect 303448 267586 303796 267618
rect 437816 268174 438164 268206
rect 437816 267938 437872 268174
rect 438108 267938 438164 268174
rect 437816 267854 438164 267938
rect 437816 267618 437872 267854
rect 438108 267618 438164 267854
rect 437816 267586 438164 267618
rect 302768 264454 303116 264486
rect 302768 264218 302824 264454
rect 303060 264218 303116 264454
rect 302768 264134 303116 264218
rect 302768 263898 302824 264134
rect 303060 263898 303116 264134
rect 302768 263866 303116 263898
rect 438496 264454 438844 264486
rect 438496 264218 438552 264454
rect 438788 264218 438844 264454
rect 438496 264134 438844 264218
rect 438496 263898 438552 264134
rect 438788 263898 438844 264134
rect 438496 263866 438844 263898
rect 441662 259317 441722 319227
rect 441659 259316 441725 259317
rect 441659 259252 441660 259316
rect 441724 259252 441725 259316
rect 441659 259251 441725 259252
rect 303448 258174 303796 258206
rect 303448 257938 303504 258174
rect 303740 257938 303796 258174
rect 303448 257854 303796 257938
rect 303448 257618 303504 257854
rect 303740 257618 303796 257854
rect 303448 257586 303796 257618
rect 437816 258174 438164 258206
rect 437816 257938 437872 258174
rect 438108 257938 438164 258174
rect 437816 257854 438164 257938
rect 437816 257618 437872 257854
rect 438108 257618 438164 257854
rect 437816 257586 438164 257618
rect 302768 254454 303116 254486
rect 302768 254218 302824 254454
rect 303060 254218 303116 254454
rect 302768 254134 303116 254218
rect 302768 253898 302824 254134
rect 303060 253898 303116 254134
rect 302768 253866 303116 253898
rect 438496 254454 438844 254486
rect 438496 254218 438552 254454
rect 438788 254218 438844 254454
rect 438496 254134 438844 254218
rect 438496 253898 438552 254134
rect 438788 253898 438844 254134
rect 438496 253866 438844 253898
rect 441659 253604 441725 253605
rect 441659 253540 441660 253604
rect 441724 253540 441725 253604
rect 441659 253539 441725 253540
rect 302371 249796 302437 249797
rect 302371 249732 302372 249796
rect 302436 249732 302437 249796
rect 302371 249731 302437 249732
rect 302003 218652 302069 218653
rect 302003 218588 302004 218652
rect 302068 218588 302069 218652
rect 302003 218587 302069 218588
rect 300531 217428 300597 217429
rect 300531 217364 300532 217428
rect 300596 217364 300597 217428
rect 300531 217363 300597 217364
rect 302374 214029 302434 249731
rect 303448 248174 303796 248206
rect 303448 247938 303504 248174
rect 303740 247938 303796 248174
rect 303448 247854 303796 247938
rect 303448 247618 303504 247854
rect 303740 247618 303796 247854
rect 303448 247586 303796 247618
rect 437816 248174 438164 248206
rect 437816 247938 437872 248174
rect 438108 247938 438164 248174
rect 437816 247854 438164 247938
rect 437816 247618 437872 247854
rect 438108 247618 438164 247854
rect 437816 247586 438164 247618
rect 302768 244454 303116 244486
rect 302768 244218 302824 244454
rect 303060 244218 303116 244454
rect 302768 244134 303116 244218
rect 302768 243898 302824 244134
rect 303060 243898 303116 244134
rect 302768 243866 303116 243898
rect 438496 244454 438844 244486
rect 438496 244218 438552 244454
rect 438788 244218 438844 244454
rect 438496 244134 438844 244218
rect 438496 243898 438552 244134
rect 438788 243898 438844 244134
rect 438496 243866 438844 243898
rect 425750 240040 425886 240070
rect 304763 240004 304829 240005
rect 304763 239940 304764 240004
rect 304828 239940 304829 240004
rect 304763 239939 304829 239940
rect 302371 214028 302437 214029
rect 302371 213964 302372 214028
rect 302436 213964 302437 214028
rect 302371 213963 302437 213964
rect 304766 212938 304826 239939
rect 318552 239730 318612 240040
rect 319640 239730 319700 240040
rect 320728 239730 320788 240040
rect 318552 239670 318626 239730
rect 319640 239670 319730 239730
rect 308259 237420 308325 237421
rect 308259 237356 308260 237420
rect 308324 237356 308325 237420
rect 308259 237355 308325 237356
rect 305683 236060 305749 236061
rect 305683 235996 305684 236060
rect 305748 235996 305749 236060
rect 305683 235995 305749 235996
rect 305131 217428 305197 217429
rect 305131 217364 305132 217428
rect 305196 217364 305197 217428
rect 305131 217363 305197 217364
rect 305134 212938 305194 217363
rect 305686 213210 305746 235995
rect 306051 229804 306117 229805
rect 306051 229740 306052 229804
rect 306116 229740 306117 229804
rect 306051 229739 306117 229740
rect 305594 213150 305746 213210
rect 304766 212878 304918 212938
rect 305134 212878 305286 212938
rect 304858 212550 304918 212878
rect 305226 212580 305286 212878
rect 304766 212490 304918 212550
rect 305134 212520 305286 212580
rect 305594 212550 305654 213150
rect 306054 212938 306114 229739
rect 307155 225044 307221 225045
rect 307155 224980 307156 225044
rect 307220 224980 307221 225044
rect 307155 224979 307221 224980
rect 306787 217292 306853 217293
rect 306787 217228 306788 217292
rect 306852 217228 306853 217292
rect 306787 217227 306853 217228
rect 306419 216068 306485 216069
rect 306419 216004 306420 216068
rect 306484 216004 306485 216068
rect 306419 216003 306485 216004
rect 306422 213210 306482 216003
rect 306790 213210 306850 217227
rect 305962 212878 306114 212938
rect 306330 213150 306482 213210
rect 306698 213150 306850 213210
rect 305962 212580 306022 212878
rect 305962 212520 306114 212580
rect 306330 212550 306390 213150
rect 306698 212550 306758 213150
rect 307158 212938 307218 224979
rect 307891 224364 307957 224365
rect 307891 224300 307892 224364
rect 307956 224300 307957 224364
rect 307891 224299 307957 224300
rect 307523 220148 307589 220149
rect 307523 220084 307524 220148
rect 307588 220084 307589 220148
rect 307523 220083 307589 220084
rect 307526 212938 307586 220083
rect 307894 212938 307954 224299
rect 308262 212938 308322 237355
rect 312491 236740 312557 236741
rect 312491 236676 312492 236740
rect 312556 236676 312557 236740
rect 312491 236675 312557 236676
rect 308995 235924 309061 235925
rect 308995 235860 308996 235924
rect 309060 235860 309061 235924
rect 308995 235859 309061 235860
rect 308998 213210 309058 235859
rect 309363 233884 309429 233885
rect 309363 233820 309364 233884
rect 309428 233820 309429 233884
rect 309363 233819 309429 233820
rect 310835 233884 310901 233885
rect 310835 233820 310836 233884
rect 310900 233820 310901 233884
rect 310835 233819 310901 233820
rect 308906 213150 309058 213210
rect 307066 212878 307218 212938
rect 307434 212878 307586 212938
rect 307802 212878 307954 212938
rect 308170 212878 308322 212938
rect 308535 212940 308601 212941
rect 307066 212580 307126 212878
rect 307066 212520 307218 212580
rect 304766 212470 304888 212490
rect 305134 212470 305256 212520
rect 305992 212470 306114 212520
rect 307096 212489 307218 212520
rect 307434 212490 307494 212878
rect 307802 212550 307862 212878
rect 308170 212550 308230 212878
rect 308535 212876 308536 212940
rect 308600 212876 308601 212940
rect 308535 212875 308601 212876
rect 307802 212490 307954 212550
rect 308170 212490 308322 212550
rect 308538 212500 308598 212875
rect 308906 212550 308966 213150
rect 309366 212938 309426 233819
rect 309731 232524 309797 232525
rect 309731 232460 309732 232524
rect 309796 232460 309797 232524
rect 309731 232459 309797 232460
rect 309734 213210 309794 232459
rect 309915 218652 309981 218653
rect 309915 218588 309916 218652
rect 309980 218588 309981 218652
rect 309915 218587 309981 218588
rect 309274 212878 309426 212938
rect 309642 213150 309794 213210
rect 309918 213210 309978 218587
rect 310283 214028 310349 214029
rect 310283 213964 310284 214028
rect 310348 213964 310349 214028
rect 310283 213963 310349 213964
rect 309918 213150 310070 213210
rect 309274 212500 309334 212878
rect 309642 212550 309702 213150
rect 310010 212550 310070 213150
rect 310286 212938 310346 213963
rect 310838 213210 310898 233819
rect 311939 225996 312005 225997
rect 311939 225932 311940 225996
rect 312004 225932 312005 225996
rect 311939 225931 312005 225932
rect 311019 222868 311085 222869
rect 311019 222804 311020 222868
rect 311084 222804 311085 222868
rect 311019 222803 311085 222804
rect 311022 216069 311082 222803
rect 311203 218652 311269 218653
rect 311203 218588 311204 218652
rect 311268 218588 311269 218652
rect 311203 218587 311269 218588
rect 311019 216068 311085 216069
rect 311019 216004 311020 216068
rect 311084 216004 311085 216068
rect 311019 216003 311085 216004
rect 310746 213150 310898 213210
rect 310286 212878 310438 212938
rect 310378 212500 310438 212878
rect 310746 212550 310806 213150
rect 311206 212938 311266 218587
rect 311942 213210 312002 225931
rect 312494 225045 312554 236675
rect 318566 236061 318626 239670
rect 316539 236060 316605 236061
rect 316539 235996 316540 236060
rect 316604 235996 316605 236060
rect 316539 235995 316605 235996
rect 318563 236060 318629 236061
rect 318563 235996 318564 236060
rect 318628 235996 318629 236060
rect 318563 235995 318629 235996
rect 319483 236060 319549 236061
rect 319483 235996 319484 236060
rect 319548 235996 319549 236060
rect 319483 235995 319549 235996
rect 313411 235516 313477 235517
rect 313411 235452 313412 235516
rect 313476 235452 313477 235516
rect 313411 235451 313477 235452
rect 312491 225044 312557 225045
rect 312491 224980 312492 225044
rect 312556 224980 312557 225044
rect 312491 224979 312557 224980
rect 312491 224228 312557 224229
rect 312491 224164 312492 224228
rect 312556 224164 312557 224228
rect 312491 224163 312557 224164
rect 312307 214572 312373 214573
rect 312307 214508 312308 214572
rect 312372 214508 312373 214572
rect 312307 214507 312373 214508
rect 311850 213150 312002 213210
rect 311479 213076 311545 213077
rect 311479 213012 311480 213076
rect 311544 213012 311545 213076
rect 311479 213011 311545 213012
rect 311114 212878 311266 212938
rect 311114 212500 311174 212878
rect 311482 212519 311542 213011
rect 311850 212550 311910 213150
rect 312310 212938 312370 214507
rect 312494 213077 312554 224163
rect 313043 221508 313109 221509
rect 313043 221444 313044 221508
rect 313108 221444 313109 221508
rect 313043 221443 313109 221444
rect 312675 215932 312741 215933
rect 312675 215868 312676 215932
rect 312740 215868 312741 215932
rect 312675 215867 312741 215868
rect 312491 213076 312557 213077
rect 312491 213012 312492 213076
rect 312556 213012 312557 213076
rect 312491 213011 312557 213012
rect 312678 212938 312738 215867
rect 313046 213210 313106 221443
rect 313414 213210 313474 235451
rect 314883 232524 314949 232525
rect 314883 232460 314884 232524
rect 314948 232460 314949 232524
rect 314883 232459 314949 232460
rect 314515 226948 314581 226949
rect 314515 226884 314516 226948
rect 314580 226884 314581 226948
rect 314515 226883 314581 226884
rect 313779 221780 313845 221781
rect 313779 221716 313780 221780
rect 313844 221716 313845 221780
rect 313779 221715 313845 221716
rect 312218 212878 312370 212938
rect 312586 212878 312738 212938
rect 312954 213150 313106 213210
rect 313322 213150 313474 213210
rect 312218 212500 312278 212878
rect 312586 212550 312646 212878
rect 312954 212550 313014 213150
rect 313322 212550 313382 213150
rect 313782 212938 313842 221715
rect 314147 216068 314213 216069
rect 314147 216004 314148 216068
rect 314212 216004 314213 216068
rect 314147 216003 314213 216004
rect 314150 212938 314210 216003
rect 314518 213210 314578 226883
rect 314886 213210 314946 232459
rect 315619 231436 315685 231437
rect 315619 231372 315620 231436
rect 315684 231372 315685 231436
rect 315619 231371 315685 231372
rect 315251 228580 315317 228581
rect 315251 228516 315252 228580
rect 315316 228516 315317 228580
rect 315251 228515 315317 228516
rect 315254 213210 315314 228515
rect 315622 213210 315682 231371
rect 315803 230076 315869 230077
rect 315803 230012 315804 230076
rect 315868 230012 315869 230076
rect 315803 230011 315869 230012
rect 313690 212878 313842 212938
rect 314058 212878 314210 212938
rect 314426 213150 314578 213210
rect 314794 213150 314946 213210
rect 315162 213150 315314 213210
rect 315530 213150 315682 213210
rect 315806 213210 315866 230011
rect 316542 220149 316602 235995
rect 318563 234020 318629 234021
rect 318563 233956 318564 234020
rect 318628 233956 318629 234020
rect 318563 233955 318629 233956
rect 317459 232796 317525 232797
rect 317459 232732 317460 232796
rect 317524 232732 317525 232796
rect 317459 232731 317525 232732
rect 317091 227220 317157 227221
rect 317091 227156 317092 227220
rect 317156 227156 317157 227220
rect 317091 227155 317157 227156
rect 316723 225724 316789 225725
rect 316723 225660 316724 225724
rect 316788 225660 316789 225724
rect 316723 225659 316789 225660
rect 316539 220148 316605 220149
rect 316539 220084 316540 220148
rect 316604 220084 316605 220148
rect 316539 220083 316605 220084
rect 316355 215252 316421 215253
rect 316355 215188 316356 215252
rect 316420 215188 316421 215252
rect 316355 215187 316421 215188
rect 315806 213150 315958 213210
rect 313690 212500 313750 212878
rect 314058 212550 314118 212878
rect 314426 212550 314486 213150
rect 314794 212550 314854 213150
rect 315162 212550 315222 213150
rect 315530 212550 315590 213150
rect 315898 212550 315958 213150
rect 316358 212938 316418 215187
rect 316726 212938 316786 225659
rect 317094 213210 317154 227155
rect 316266 212878 316418 212938
rect 316634 212878 316786 212938
rect 317002 213150 317154 213210
rect 316266 212500 316326 212878
rect 316634 212500 316694 212878
rect 317002 212550 317062 213150
rect 317462 213074 317522 232731
rect 318195 231300 318261 231301
rect 318195 231236 318196 231300
rect 318260 231236 318261 231300
rect 318195 231235 318261 231236
rect 317827 228308 317893 228309
rect 317827 228244 317828 228308
rect 317892 228244 317893 228308
rect 317827 228243 317893 228244
rect 317830 213210 317890 228243
rect 318198 213210 318258 231235
rect 318566 213210 318626 233955
rect 318931 217564 318997 217565
rect 318931 217500 318932 217564
rect 318996 217500 318997 217564
rect 318931 217499 318997 217500
rect 318934 213210 318994 217499
rect 319299 217428 319365 217429
rect 319299 217364 319300 217428
rect 319364 217364 319365 217428
rect 319299 217363 319365 217364
rect 317370 213014 317522 213074
rect 317738 213150 317890 213210
rect 318106 213150 318258 213210
rect 318474 213150 318626 213210
rect 318842 213150 318994 213210
rect 317370 212500 317430 213014
rect 317738 212550 317798 213150
rect 318106 212550 318166 213150
rect 318474 212550 318534 213150
rect 318842 212550 318902 213150
rect 319302 213074 319362 217363
rect 319486 217293 319546 235995
rect 319670 224365 319730 239670
rect 320590 239670 320788 239730
rect 322088 239730 322148 240040
rect 323040 239730 323100 240040
rect 322088 239670 322306 239730
rect 320590 229805 320650 239670
rect 320771 235244 320837 235245
rect 320771 235180 320772 235244
rect 320836 235180 320837 235244
rect 320771 235179 320837 235180
rect 320587 229804 320653 229805
rect 320587 229740 320588 229804
rect 320652 229740 320653 229804
rect 320587 229739 320653 229740
rect 319667 224364 319733 224365
rect 319667 224300 319668 224364
rect 319732 224300 319733 224364
rect 319667 224299 319733 224300
rect 320035 220420 320101 220421
rect 320035 220356 320036 220420
rect 320100 220356 320101 220420
rect 320035 220355 320101 220356
rect 319667 218788 319733 218789
rect 319667 218724 319668 218788
rect 319732 218724 319733 218788
rect 319667 218723 319733 218724
rect 319483 217292 319549 217293
rect 319483 217228 319484 217292
rect 319548 217228 319549 217292
rect 319483 217227 319549 217228
rect 319210 213014 319362 213074
rect 319210 212500 319270 213014
rect 319670 212938 319730 218723
rect 320038 213074 320098 220355
rect 320403 220284 320469 220285
rect 320403 220220 320404 220284
rect 320468 220220 320469 220284
rect 320403 220219 320469 220220
rect 319578 212878 319730 212938
rect 319946 213014 320098 213074
rect 319578 212550 319638 212878
rect 319946 212500 320006 213014
rect 320406 212938 320466 220219
rect 320774 213210 320834 235179
rect 321875 232660 321941 232661
rect 321875 232596 321876 232660
rect 321940 232596 321941 232660
rect 321875 232595 321941 232596
rect 321139 229940 321205 229941
rect 321139 229876 321140 229940
rect 321204 229876 321205 229940
rect 321139 229875 321205 229876
rect 321142 213210 321202 229875
rect 321323 227084 321389 227085
rect 321323 227020 321324 227084
rect 321388 227020 321389 227084
rect 321323 227019 321389 227020
rect 320314 212878 320466 212938
rect 320682 213150 320834 213210
rect 321050 213150 321202 213210
rect 321326 213210 321386 227019
rect 321878 213210 321938 232595
rect 322246 222869 322306 239670
rect 322982 239670 323100 239730
rect 324264 239730 324324 240040
rect 325624 239730 325684 240040
rect 324264 239670 324330 239730
rect 322982 236061 323042 239670
rect 324270 236741 324330 239670
rect 325558 239670 325684 239730
rect 326712 239730 326772 240040
rect 327936 239730 327996 240040
rect 329024 239730 329084 240040
rect 330112 239730 330172 240040
rect 330792 239730 330852 240040
rect 331200 239730 331260 240040
rect 332560 239730 332620 240040
rect 333240 239730 333300 240040
rect 333784 239730 333844 240040
rect 334872 239730 334932 240040
rect 335960 239730 336020 240040
rect 326712 239670 326906 239730
rect 327936 239670 328010 239730
rect 329024 239670 329114 239730
rect 330112 239670 330218 239730
rect 330792 239670 330954 239730
rect 331200 239670 331322 239730
rect 332560 239670 332794 239730
rect 333240 239670 333346 239730
rect 333784 239670 333898 239730
rect 334872 239670 335002 239730
rect 324267 236740 324333 236741
rect 324267 236676 324268 236740
rect 324332 236676 324333 236740
rect 324267 236675 324333 236676
rect 325371 236740 325437 236741
rect 325371 236676 325372 236740
rect 325436 236676 325437 236740
rect 325371 236675 325437 236676
rect 323531 236604 323597 236605
rect 323531 236540 323532 236604
rect 323596 236540 323597 236604
rect 323531 236539 323597 236540
rect 322979 236060 323045 236061
rect 322979 235996 322980 236060
rect 323044 235996 323045 236060
rect 322979 235995 323045 235996
rect 323163 236060 323229 236061
rect 323163 235996 323164 236060
rect 323228 235996 323229 236060
rect 323163 235995 323229 235996
rect 323166 233885 323226 235995
rect 323163 233884 323229 233885
rect 323163 233820 323164 233884
rect 323228 233820 323229 233884
rect 323163 233819 323229 233820
rect 323534 226949 323594 236539
rect 323715 235652 323781 235653
rect 323715 235588 323716 235652
rect 323780 235588 323781 235652
rect 323715 235587 323781 235588
rect 323531 226948 323597 226949
rect 323531 226884 323532 226948
rect 323596 226884 323597 226948
rect 323531 226883 323597 226884
rect 322611 223276 322677 223277
rect 322611 223212 322612 223276
rect 322676 223212 322677 223276
rect 322611 223211 322677 223212
rect 322243 222868 322309 222869
rect 322243 222804 322244 222868
rect 322308 222804 322309 222868
rect 322243 222803 322309 222804
rect 322243 221644 322309 221645
rect 322243 221580 322244 221644
rect 322308 221580 322309 221644
rect 322243 221579 322309 221580
rect 322246 213210 322306 221579
rect 321326 213150 321478 213210
rect 320314 212550 320374 212878
rect 320682 212550 320742 213150
rect 321050 212550 321110 213150
rect 321418 212550 321478 213150
rect 321786 213150 321938 213210
rect 322154 213150 322306 213210
rect 321786 212550 321846 213150
rect 322154 212550 322214 213150
rect 322614 213074 322674 223211
rect 323347 223004 323413 223005
rect 323347 222940 323348 223004
rect 323412 222940 323413 223004
rect 323347 222939 323413 222940
rect 323350 213210 323410 222939
rect 323258 213150 323410 213210
rect 322522 213014 322674 213074
rect 322887 213076 322953 213077
rect 322522 212500 322582 213014
rect 322887 213012 322888 213076
rect 322952 213012 322953 213076
rect 322887 213011 322953 213012
rect 322890 212550 322950 213011
rect 323258 212550 323318 213150
rect 323718 213074 323778 235587
rect 325003 234156 325069 234157
rect 325003 234092 325004 234156
rect 325068 234092 325069 234156
rect 325003 234091 325069 234092
rect 324819 225860 324885 225861
rect 324819 225796 324820 225860
rect 324884 225796 324885 225860
rect 324819 225795 324885 225796
rect 324083 224500 324149 224501
rect 324083 224436 324084 224500
rect 324148 224436 324149 224500
rect 324083 224435 324149 224436
rect 324086 213074 324146 224435
rect 324267 219060 324333 219061
rect 324267 218996 324268 219060
rect 324332 218996 324333 219060
rect 324267 218995 324333 218996
rect 324270 216069 324330 218995
rect 324451 216204 324517 216205
rect 324451 216140 324452 216204
rect 324516 216140 324517 216204
rect 324451 216139 324517 216140
rect 324267 216068 324333 216069
rect 324267 216004 324268 216068
rect 324332 216004 324333 216068
rect 324267 216003 324333 216004
rect 323626 213014 323778 213074
rect 323994 213014 324146 213074
rect 323626 212500 323686 213014
rect 323994 212500 324054 213014
rect 324454 212938 324514 216139
rect 324822 213210 324882 225795
rect 325006 215253 325066 234091
rect 325374 229110 325434 236675
rect 325558 236061 325618 239670
rect 325555 236060 325621 236061
rect 325555 235996 325556 236060
rect 325620 235996 325621 236060
rect 325555 235995 325621 235996
rect 326659 231164 326725 231165
rect 326659 231100 326660 231164
rect 326724 231100 326725 231164
rect 326659 231099 326725 231100
rect 326475 230484 326541 230485
rect 326475 230420 326476 230484
rect 326540 230420 326541 230484
rect 326475 230419 326541 230420
rect 325374 229050 325618 229110
rect 325003 215252 325069 215253
rect 325003 215188 325004 215252
rect 325068 215188 325069 215252
rect 325003 215187 325069 215188
rect 325187 214844 325253 214845
rect 325187 214780 325188 214844
rect 325252 214780 325253 214844
rect 325187 214779 325253 214780
rect 324362 212878 324514 212938
rect 324730 213150 324882 213210
rect 324362 212550 324422 212878
rect 324730 212550 324790 213150
rect 325190 213074 325250 214779
rect 325558 213210 325618 229050
rect 325923 216748 325989 216749
rect 325923 216684 325924 216748
rect 325988 216684 325989 216748
rect 325923 216683 325989 216684
rect 325098 213014 325250 213074
rect 325466 213150 325618 213210
rect 325098 212500 325158 213014
rect 325466 212550 325526 213150
rect 325926 212938 325986 216683
rect 326478 213213 326538 230419
rect 326662 222210 326722 231099
rect 326846 229110 326906 239670
rect 327395 233884 327461 233885
rect 327395 233820 327396 233884
rect 327460 233820 327461 233884
rect 327395 233819 327461 233820
rect 326846 229050 327090 229110
rect 326662 222150 326906 222210
rect 326659 218924 326725 218925
rect 326659 218860 326660 218924
rect 326724 218860 326725 218924
rect 326659 218859 326725 218860
rect 326475 213212 326541 213213
rect 326475 213148 326476 213212
rect 326540 213148 326541 213212
rect 326475 213147 326541 213148
rect 326199 213076 326265 213077
rect 326199 213012 326200 213076
rect 326264 213012 326265 213076
rect 326199 213011 326265 213012
rect 325834 212878 325986 212938
rect 325834 212550 325894 212878
rect 326202 212550 326262 213011
rect 326662 212938 326722 218859
rect 326846 213210 326906 222150
rect 327030 218653 327090 229050
rect 327027 218652 327093 218653
rect 327027 218588 327028 218652
rect 327092 218588 327093 218652
rect 327027 218587 327093 218588
rect 326846 213150 326998 213210
rect 326570 212878 326722 212938
rect 326570 212500 326630 212878
rect 326938 212550 326998 213150
rect 327398 213074 327458 233819
rect 327579 228444 327645 228445
rect 327579 228380 327580 228444
rect 327644 228380 327645 228444
rect 327579 228379 327645 228380
rect 327582 213077 327642 228379
rect 327950 224229 328010 239670
rect 329054 225997 329114 239670
rect 329419 236876 329485 236877
rect 329419 236812 329420 236876
rect 329484 236812 329485 236876
rect 329419 236811 329485 236812
rect 329051 225996 329117 225997
rect 329051 225932 329052 225996
rect 329116 225932 329117 225996
rect 329051 225931 329117 225932
rect 328499 225588 328565 225589
rect 328499 225524 328500 225588
rect 328564 225524 328565 225588
rect 328499 225523 328565 225524
rect 327947 224228 328013 224229
rect 327947 224164 327948 224228
rect 328012 224164 328013 224228
rect 327947 224163 328013 224164
rect 328315 224228 328381 224229
rect 328315 224164 328316 224228
rect 328380 224164 328381 224228
rect 328315 224163 328381 224164
rect 328318 216069 328378 224163
rect 328315 216068 328381 216069
rect 328315 216004 328316 216068
rect 328380 216004 328381 216068
rect 328315 216003 328381 216004
rect 328502 215930 328562 225523
rect 329235 220148 329301 220149
rect 329235 220084 329236 220148
rect 329300 220084 329301 220148
rect 329235 220083 329301 220084
rect 328683 216068 328749 216069
rect 328683 216004 328684 216068
rect 328748 216004 328749 216068
rect 328683 216003 328749 216004
rect 328134 215870 328562 215930
rect 328134 213210 328194 215870
rect 328686 213210 328746 216003
rect 329238 213210 329298 220083
rect 329422 216749 329482 236811
rect 329603 217292 329669 217293
rect 329603 217228 329604 217292
rect 329668 217228 329669 217292
rect 329603 217227 329669 217228
rect 329419 216748 329485 216749
rect 329419 216684 329420 216748
rect 329484 216684 329485 216748
rect 329419 216683 329485 216684
rect 329606 213210 329666 217227
rect 329971 215932 330037 215933
rect 329971 215868 329972 215932
rect 330036 215868 330037 215932
rect 329971 215867 330037 215868
rect 329974 213210 330034 215867
rect 330158 214573 330218 239670
rect 330894 223277 330954 239670
rect 331262 224229 331322 239670
rect 331995 226948 332061 226949
rect 331995 226884 331996 226948
rect 332060 226884 332061 226948
rect 331995 226883 332061 226884
rect 331443 224364 331509 224365
rect 331443 224300 331444 224364
rect 331508 224300 331509 224364
rect 331443 224299 331509 224300
rect 331259 224228 331325 224229
rect 331259 224164 331260 224228
rect 331324 224164 331325 224228
rect 331259 224163 331325 224164
rect 330891 223276 330957 223277
rect 330891 223212 330892 223276
rect 330956 223212 330957 223276
rect 330891 223211 330957 223212
rect 330523 223140 330589 223141
rect 330523 223076 330524 223140
rect 330588 223076 330589 223140
rect 330523 223075 330589 223076
rect 330339 222868 330405 222869
rect 330339 222804 330340 222868
rect 330404 222804 330405 222868
rect 330339 222803 330405 222804
rect 330155 214572 330221 214573
rect 330155 214508 330156 214572
rect 330220 214508 330221 214572
rect 330155 214507 330221 214508
rect 330342 213210 330402 222803
rect 330526 216205 330586 223075
rect 331075 218652 331141 218653
rect 331075 218588 331076 218652
rect 331140 218588 331141 218652
rect 331075 218587 331141 218588
rect 330707 217156 330773 217157
rect 330707 217092 330708 217156
rect 330772 217092 330773 217156
rect 330707 217091 330773 217092
rect 330523 216204 330589 216205
rect 330523 216140 330524 216204
rect 330588 216140 330589 216204
rect 330523 216139 330589 216140
rect 330710 213210 330770 217091
rect 331078 213210 331138 218587
rect 331446 213210 331506 224299
rect 331998 217157 332058 226883
rect 332363 224228 332429 224229
rect 332363 224164 332364 224228
rect 332428 224164 332429 224228
rect 332363 224163 332429 224164
rect 331995 217156 332061 217157
rect 331995 217092 331996 217156
rect 332060 217092 332061 217156
rect 331995 217091 332061 217092
rect 332179 214708 332245 214709
rect 332179 214644 332180 214708
rect 332244 214644 332245 214708
rect 332179 214643 332245 214644
rect 331811 214572 331877 214573
rect 331811 214508 331812 214572
rect 331876 214508 331877 214572
rect 331811 214507 331877 214508
rect 331814 213210 331874 214507
rect 332182 213210 332242 214643
rect 328042 213150 328194 213210
rect 328410 213150 328746 213210
rect 329146 213150 329298 213210
rect 329514 213150 329666 213210
rect 329882 213150 330034 213210
rect 330250 213150 330402 213210
rect 330618 213150 330770 213210
rect 330986 213150 331138 213210
rect 331354 213150 331506 213210
rect 331722 213150 331874 213210
rect 332090 213150 332242 213210
rect 332366 213210 332426 224163
rect 332734 221509 332794 239670
rect 333099 235380 333165 235381
rect 333099 235316 333100 235380
rect 333164 235316 333165 235380
rect 333099 235315 333165 235316
rect 332731 221508 332797 221509
rect 332731 221444 332732 221508
rect 332796 221444 332797 221508
rect 332731 221443 332797 221444
rect 332915 216204 332981 216205
rect 332915 216140 332916 216204
rect 332980 216140 332981 216204
rect 332915 216139 332981 216140
rect 332918 213210 332978 216139
rect 333102 215797 333162 235315
rect 333286 230485 333346 239670
rect 333838 235517 333898 239670
rect 334571 236060 334637 236061
rect 334571 235996 334572 236060
rect 334636 235996 334637 236060
rect 334571 235995 334637 235996
rect 333835 235516 333901 235517
rect 333835 235452 333836 235516
rect 333900 235452 333901 235516
rect 333835 235451 333901 235452
rect 333283 230484 333349 230485
rect 333283 230420 333284 230484
rect 333348 230420 333349 230484
rect 333283 230419 333349 230420
rect 333651 229804 333717 229805
rect 333651 229740 333652 229804
rect 333716 229740 333717 229804
rect 333651 229739 333717 229740
rect 333283 221508 333349 221509
rect 333283 221444 333284 221508
rect 333348 221444 333349 221508
rect 333283 221443 333349 221444
rect 333099 215796 333165 215797
rect 333099 215732 333100 215796
rect 333164 215732 333165 215796
rect 333099 215731 333165 215732
rect 333286 213210 333346 221443
rect 333654 213210 333714 229739
rect 334574 223005 334634 235995
rect 334571 223004 334637 223005
rect 334571 222940 334572 223004
rect 334636 222940 334637 223004
rect 334571 222939 334637 222940
rect 334755 223004 334821 223005
rect 334755 222940 334756 223004
rect 334820 222940 334821 223004
rect 334755 222939 334821 222940
rect 334571 221916 334637 221917
rect 334571 221852 334572 221916
rect 334636 221852 334637 221916
rect 334571 221851 334637 221852
rect 332366 213150 332518 213210
rect 327306 213014 327458 213074
rect 327579 213076 327645 213077
rect 327306 212500 327366 213014
rect 327579 213012 327580 213076
rect 327644 213012 327645 213076
rect 327579 213011 327645 213012
rect 327671 212940 327737 212941
rect 327671 212876 327672 212940
rect 327736 212876 327737 212940
rect 327671 212875 327737 212876
rect 327674 212550 327734 212875
rect 328042 212550 328102 213150
rect 328410 212550 328470 213150
rect 328775 213076 328841 213077
rect 328775 213012 328776 213076
rect 328840 213012 328841 213076
rect 328775 213011 328841 213012
rect 328778 212500 328838 213011
rect 329146 212550 329206 213150
rect 329514 212550 329574 213150
rect 329882 212550 329942 213150
rect 330250 212550 330310 213150
rect 330618 212550 330678 213150
rect 330986 212550 331046 213150
rect 331354 212550 331414 213150
rect 329146 212490 329298 212550
rect 329514 212490 329666 212550
rect 330250 212490 330402 212550
rect 330618 212490 330770 212550
rect 331722 212490 331782 213150
rect 332090 212490 332150 213150
rect 332458 212550 332518 213150
rect 332826 213150 332978 213210
rect 333194 213150 333346 213210
rect 333562 213150 333714 213210
rect 332826 212550 332886 213150
rect 333194 212550 333254 213150
rect 333562 212550 333622 213150
rect 334574 212580 334634 221851
rect 334758 213077 334818 222939
rect 334942 221781 335002 239670
rect 335862 239670 336020 239730
rect 336096 239730 336156 240040
rect 337048 239730 337108 240040
rect 338408 239730 338468 240040
rect 336096 239670 336290 239730
rect 335862 238770 335922 239670
rect 335862 238710 336106 238770
rect 334939 221780 335005 221781
rect 334939 221716 334940 221780
rect 335004 221716 335005 221780
rect 334939 221715 335005 221716
rect 336046 219061 336106 238710
rect 336230 236061 336290 239670
rect 336966 239670 337108 239730
rect 338254 239670 338468 239730
rect 338544 239730 338604 240040
rect 339496 239730 339556 240040
rect 340584 239730 340644 240040
rect 338544 239670 338682 239730
rect 339496 239670 339602 239730
rect 336966 236605 337026 239670
rect 337331 237964 337397 237965
rect 337331 237900 337332 237964
rect 337396 237900 337397 237964
rect 337331 237899 337397 237900
rect 336963 236604 337029 236605
rect 336963 236540 336964 236604
rect 337028 236540 337029 236604
rect 336963 236539 337029 236540
rect 336227 236060 336293 236061
rect 336227 235996 336228 236060
rect 336292 235996 336293 236060
rect 336227 235995 336293 235996
rect 336043 219060 336109 219061
rect 336043 218996 336044 219060
rect 336108 218996 336109 219060
rect 336043 218995 336109 218996
rect 334755 213076 334821 213077
rect 334755 213012 334756 213076
rect 334820 213012 334821 213076
rect 334755 213011 334821 213012
rect 333960 212520 334634 212580
rect 307832 212470 307954 212490
rect 308200 212470 308322 212490
rect 329176 212470 329298 212490
rect 329544 212470 329666 212490
rect 330280 212470 330402 212490
rect 330648 212470 330770 212490
rect 307365 208174 307685 208206
rect 307365 207938 307407 208174
rect 307643 207938 307685 208174
rect 307365 207854 307685 207938
rect 307365 207618 307407 207854
rect 307643 207618 307685 207854
rect 307365 207586 307685 207618
rect 315207 208174 315527 208206
rect 315207 207938 315249 208174
rect 315485 207938 315527 208174
rect 315207 207854 315527 207938
rect 315207 207618 315249 207854
rect 315485 207618 315527 207854
rect 315207 207586 315527 207618
rect 323049 208174 323369 208206
rect 323049 207938 323091 208174
rect 323327 207938 323369 208174
rect 323049 207854 323369 207938
rect 323049 207618 323091 207854
rect 323327 207618 323369 207854
rect 323049 207586 323369 207618
rect 330891 208174 331211 208206
rect 330891 207938 330933 208174
rect 331169 207938 331211 208174
rect 330891 207854 331211 207938
rect 330891 207618 330933 207854
rect 331169 207618 331211 207854
rect 330891 207586 331211 207618
rect 303444 204454 303764 204486
rect 303444 204218 303486 204454
rect 303722 204218 303764 204454
rect 303444 204134 303764 204218
rect 303444 203898 303486 204134
rect 303722 203898 303764 204134
rect 303444 203866 303764 203898
rect 311286 204454 311606 204486
rect 311286 204218 311328 204454
rect 311564 204218 311606 204454
rect 311286 204134 311606 204218
rect 311286 203898 311328 204134
rect 311564 203898 311606 204134
rect 311286 203866 311606 203898
rect 319128 204454 319448 204486
rect 319128 204218 319170 204454
rect 319406 204218 319448 204454
rect 319128 204134 319448 204218
rect 319128 203898 319170 204134
rect 319406 203898 319448 204134
rect 319128 203866 319448 203898
rect 326970 204454 327290 204486
rect 326970 204218 327012 204454
rect 327248 204218 327290 204454
rect 326970 204134 327290 204218
rect 326970 203898 327012 204134
rect 327248 203898 327290 204134
rect 326970 203866 327290 203898
rect 307365 198174 307685 198206
rect 307365 197938 307407 198174
rect 307643 197938 307685 198174
rect 307365 197854 307685 197938
rect 307365 197618 307407 197854
rect 307643 197618 307685 197854
rect 307365 197586 307685 197618
rect 315207 198174 315527 198206
rect 315207 197938 315249 198174
rect 315485 197938 315527 198174
rect 315207 197854 315527 197938
rect 315207 197618 315249 197854
rect 315485 197618 315527 197854
rect 315207 197586 315527 197618
rect 323049 198174 323369 198206
rect 323049 197938 323091 198174
rect 323327 197938 323369 198174
rect 323049 197854 323369 197938
rect 323049 197618 323091 197854
rect 323327 197618 323369 197854
rect 323049 197586 323369 197618
rect 330891 198174 331211 198206
rect 330891 197938 330933 198174
rect 331169 197938 331211 198174
rect 330891 197854 331211 197938
rect 330891 197618 330933 197854
rect 331169 197618 331211 197854
rect 330891 197586 331211 197618
rect 303444 194454 303764 194486
rect 303444 194218 303486 194454
rect 303722 194218 303764 194454
rect 303444 194134 303764 194218
rect 303444 193898 303486 194134
rect 303722 193898 303764 194134
rect 303444 193866 303764 193898
rect 311286 194454 311606 194486
rect 311286 194218 311328 194454
rect 311564 194218 311606 194454
rect 311286 194134 311606 194218
rect 311286 193898 311328 194134
rect 311564 193898 311606 194134
rect 311286 193866 311606 193898
rect 319128 194454 319448 194486
rect 319128 194218 319170 194454
rect 319406 194218 319448 194454
rect 319128 194134 319448 194218
rect 319128 193898 319170 194134
rect 319406 193898 319448 194134
rect 319128 193866 319448 193898
rect 326970 194454 327290 194486
rect 326970 194218 327012 194454
rect 327248 194218 327290 194454
rect 326970 194134 327290 194218
rect 326970 193898 327012 194134
rect 327248 193898 327290 194134
rect 326970 193866 327290 193898
rect 337334 191861 337394 237899
rect 337883 236196 337949 236197
rect 337883 236132 337884 236196
rect 337948 236132 337949 236196
rect 337883 236131 337949 236132
rect 337886 231437 337946 236131
rect 338254 232525 338314 239670
rect 338622 235653 338682 239670
rect 338619 235652 338685 235653
rect 338619 235588 338620 235652
rect 338684 235588 338685 235652
rect 338619 235587 338685 235588
rect 338251 232524 338317 232525
rect 338251 232460 338252 232524
rect 338316 232460 338317 232524
rect 338251 232459 338317 232460
rect 338619 232524 338685 232525
rect 338619 232460 338620 232524
rect 338684 232460 338685 232524
rect 338619 232459 338685 232460
rect 337883 231436 337949 231437
rect 337883 231372 337884 231436
rect 337948 231372 337949 231436
rect 337883 231371 337949 231372
rect 338622 216205 338682 232459
rect 339542 228581 339602 239670
rect 340462 239670 340644 239730
rect 340992 239730 341052 240040
rect 341944 239730 342004 240040
rect 343168 239730 343228 240040
rect 343576 239730 343636 240040
rect 344256 239730 344316 240040
rect 340992 239670 341074 239730
rect 341944 239670 342178 239730
rect 343168 239670 343282 239730
rect 343576 239670 343650 239730
rect 340462 236197 340522 239670
rect 340459 236196 340525 236197
rect 340459 236132 340460 236196
rect 340524 236132 340525 236196
rect 340459 236131 340525 236132
rect 340275 236060 340341 236061
rect 340275 235996 340276 236060
rect 340340 235996 340341 236060
rect 340275 235995 340341 235996
rect 339539 228580 339605 228581
rect 339539 228516 339540 228580
rect 339604 228516 339605 228580
rect 339539 228515 339605 228516
rect 340091 225996 340157 225997
rect 340091 225932 340092 225996
rect 340156 225932 340157 225996
rect 340091 225931 340157 225932
rect 338619 216204 338685 216205
rect 338619 216140 338620 216204
rect 338684 216140 338685 216204
rect 338619 216139 338685 216140
rect 340094 214845 340154 225931
rect 340278 225725 340338 235995
rect 340275 225724 340341 225725
rect 340275 225660 340276 225724
rect 340340 225660 340341 225724
rect 340275 225659 340341 225660
rect 341014 224501 341074 239670
rect 342118 230077 342178 239670
rect 343222 234157 343282 239670
rect 343219 234156 343285 234157
rect 343219 234092 343220 234156
rect 343284 234092 343285 234156
rect 343219 234091 343285 234092
rect 342115 230076 342181 230077
rect 342115 230012 342116 230076
rect 342180 230012 342181 230076
rect 342115 230011 342181 230012
rect 341011 224500 341077 224501
rect 341011 224436 341012 224500
rect 341076 224436 341077 224500
rect 341011 224435 341077 224436
rect 343590 223141 343650 239670
rect 344142 239670 344316 239730
rect 345344 239730 345404 240040
rect 346024 239730 346084 240040
rect 346432 239730 346492 240040
rect 345344 239670 345490 239730
rect 346024 239670 346226 239730
rect 344142 236061 344202 239670
rect 344139 236060 344205 236061
rect 344139 235996 344140 236060
rect 344204 235996 344205 236060
rect 344139 235995 344205 235996
rect 345430 227221 345490 239670
rect 345427 227220 345493 227221
rect 345427 227156 345428 227220
rect 345492 227156 345493 227220
rect 345427 227155 345493 227156
rect 346166 225861 346226 239670
rect 346350 239670 346492 239730
rect 347792 239730 347852 240040
rect 348472 239730 348532 240040
rect 348880 239730 348940 240040
rect 350104 239730 350164 240040
rect 350784 239730 350844 240040
rect 347792 239670 347882 239730
rect 348472 239670 348618 239730
rect 348880 239670 348986 239730
rect 346350 232797 346410 239670
rect 346347 232796 346413 232797
rect 346347 232732 346348 232796
rect 346412 232732 346413 232796
rect 346347 232731 346413 232732
rect 347822 228309 347882 239670
rect 347819 228308 347885 228309
rect 347819 228244 347820 228308
rect 347884 228244 347885 228308
rect 347819 228243 347885 228244
rect 348558 225997 348618 239670
rect 348926 231301 348986 239670
rect 350030 239670 350164 239730
rect 350766 239670 350844 239730
rect 351192 239730 351252 240040
rect 352280 239730 352340 240040
rect 353504 239730 353564 240040
rect 351192 239670 351378 239730
rect 352280 239670 352482 239730
rect 349659 236604 349725 236605
rect 349659 236540 349660 236604
rect 349724 236540 349725 236604
rect 349659 236539 349725 236540
rect 348923 231300 348989 231301
rect 348923 231236 348924 231300
rect 348988 231236 348989 231300
rect 348923 231235 348989 231236
rect 348555 225996 348621 225997
rect 348555 225932 348556 225996
rect 348620 225932 348621 225996
rect 348555 225931 348621 225932
rect 346163 225860 346229 225861
rect 346163 225796 346164 225860
rect 346228 225796 346229 225860
rect 346163 225795 346229 225796
rect 343587 223140 343653 223141
rect 343587 223076 343588 223140
rect 343652 223076 343653 223140
rect 343587 223075 343653 223076
rect 349662 221917 349722 236539
rect 350030 234021 350090 239670
rect 350766 236741 350826 239670
rect 350763 236740 350829 236741
rect 350763 236676 350764 236740
rect 350828 236676 350829 236740
rect 350763 236675 350829 236676
rect 350027 234020 350093 234021
rect 350027 233956 350028 234020
rect 350092 233956 350093 234020
rect 350027 233955 350093 233956
rect 349659 221916 349725 221917
rect 349659 221852 349660 221916
rect 349724 221852 349725 221916
rect 349659 221851 349725 221852
rect 351318 217565 351378 239670
rect 351315 217564 351381 217565
rect 351315 217500 351316 217564
rect 351380 217500 351381 217564
rect 351315 217499 351381 217500
rect 352422 217429 352482 239670
rect 353342 239670 353564 239730
rect 353640 239730 353700 240040
rect 354728 239730 354788 240040
rect 353640 239670 353770 239730
rect 353342 236877 353402 239670
rect 353339 236876 353405 236877
rect 353339 236812 353340 236876
rect 353404 236812 353405 236876
rect 353339 236811 353405 236812
rect 353710 218789 353770 239670
rect 354446 239670 354788 239730
rect 355816 239730 355876 240040
rect 356088 239730 356148 240040
rect 356904 239730 356964 240040
rect 355816 239670 355978 239730
rect 356088 239670 356162 239730
rect 354446 220421 354506 239670
rect 354443 220420 354509 220421
rect 354443 220356 354444 220420
rect 354508 220356 354509 220420
rect 354443 220355 354509 220356
rect 355918 220285 355978 239670
rect 356102 228445 356162 239670
rect 356838 239670 356964 239730
rect 358264 239730 358324 240040
rect 358536 239730 358596 240040
rect 359488 239730 359548 240040
rect 360576 239730 360636 240040
rect 358264 239670 358370 239730
rect 358536 239670 358738 239730
rect 359488 239670 359658 239730
rect 356838 235245 356898 239670
rect 356835 235244 356901 235245
rect 356835 235180 356836 235244
rect 356900 235180 356901 235244
rect 356835 235179 356901 235180
rect 358310 229941 358370 239670
rect 358307 229940 358373 229941
rect 358307 229876 358308 229940
rect 358372 229876 358373 229940
rect 358307 229875 358373 229876
rect 356099 228444 356165 228445
rect 356099 228380 356100 228444
rect 356164 228380 356165 228444
rect 356099 228379 356165 228380
rect 356651 228308 356717 228309
rect 356651 228244 356652 228308
rect 356716 228244 356717 228308
rect 356651 228243 356717 228244
rect 355915 220284 355981 220285
rect 355915 220220 355916 220284
rect 355980 220220 355981 220284
rect 355915 220219 355981 220220
rect 353707 218788 353773 218789
rect 353707 218724 353708 218788
rect 353772 218724 353773 218788
rect 353707 218723 353773 218724
rect 352419 217428 352485 217429
rect 352419 217364 352420 217428
rect 352484 217364 352485 217428
rect 352419 217363 352485 217364
rect 340091 214844 340157 214845
rect 340091 214780 340092 214844
rect 340156 214780 340157 214844
rect 340091 214779 340157 214780
rect 356654 214709 356714 228243
rect 358678 218925 358738 239670
rect 359598 227085 359658 239670
rect 360518 239670 360636 239730
rect 360984 239730 361044 240040
rect 361664 239730 361724 240040
rect 363432 239730 363492 240040
rect 366016 239730 366076 240040
rect 368464 239730 368524 240040
rect 370776 239730 370836 240040
rect 373496 239730 373556 240040
rect 375944 239730 376004 240040
rect 378392 239730 378452 240040
rect 380976 239730 381036 240040
rect 383424 239730 383484 240040
rect 386008 239730 386068 240040
rect 388456 239730 388516 240040
rect 391040 239730 391100 240040
rect 393488 239730 393548 240040
rect 395936 239730 395996 240040
rect 360984 239670 361130 239730
rect 361664 239670 361866 239730
rect 363432 239670 363522 239730
rect 366016 239670 366098 239730
rect 368464 239670 368674 239730
rect 370776 239670 370882 239730
rect 373496 239670 373642 239730
rect 375944 239670 376034 239730
rect 378392 239670 378610 239730
rect 380976 239670 381186 239730
rect 383424 239670 383578 239730
rect 386008 239670 386154 239730
rect 388456 239670 388546 239730
rect 391040 239670 391122 239730
rect 393488 239670 393698 239730
rect 360518 232661 360578 239670
rect 360515 232660 360581 232661
rect 360515 232596 360516 232660
rect 360580 232596 360581 232660
rect 360515 232595 360581 232596
rect 360699 231300 360765 231301
rect 360699 231236 360700 231300
rect 360764 231236 360765 231300
rect 360699 231235 360765 231236
rect 359595 227084 359661 227085
rect 359595 227020 359596 227084
rect 359660 227020 359661 227084
rect 359595 227019 359661 227020
rect 358675 218924 358741 218925
rect 358675 218860 358676 218924
rect 358740 218860 358741 218924
rect 358675 218859 358741 218860
rect 360702 216069 360762 231235
rect 361070 231165 361130 239670
rect 361067 231164 361133 231165
rect 361067 231100 361068 231164
rect 361132 231100 361133 231164
rect 361067 231099 361133 231100
rect 361806 221645 361866 239670
rect 363462 233885 363522 239670
rect 366038 235381 366098 239670
rect 366035 235380 366101 235381
rect 366035 235316 366036 235380
rect 366100 235316 366101 235380
rect 366035 235315 366101 235316
rect 363459 233884 363525 233885
rect 363459 233820 363460 233884
rect 363524 233820 363525 233884
rect 363459 233819 363525 233820
rect 368614 225589 368674 239670
rect 370822 231301 370882 239670
rect 370819 231300 370885 231301
rect 370819 231236 370820 231300
rect 370884 231236 370885 231300
rect 370819 231235 370885 231236
rect 368611 225588 368677 225589
rect 368611 225524 368612 225588
rect 368676 225524 368677 225588
rect 368611 225523 368677 225524
rect 373582 223005 373642 239670
rect 373579 223004 373645 223005
rect 373579 222940 373580 223004
rect 373644 222940 373645 223004
rect 373579 222939 373645 222940
rect 361803 221644 361869 221645
rect 361803 221580 361804 221644
rect 361868 221580 361869 221644
rect 361803 221579 361869 221580
rect 375974 220149 376034 239670
rect 375971 220148 376037 220149
rect 375971 220084 375972 220148
rect 376036 220084 376037 220148
rect 375971 220083 376037 220084
rect 378550 217293 378610 239670
rect 378547 217292 378613 217293
rect 378547 217228 378548 217292
rect 378612 217228 378613 217292
rect 378547 217227 378613 217228
rect 360699 216068 360765 216069
rect 360699 216004 360700 216068
rect 360764 216004 360765 216068
rect 360699 216003 360765 216004
rect 381126 215933 381186 239670
rect 383518 222869 383578 239670
rect 386094 226949 386154 239670
rect 386091 226948 386157 226949
rect 386091 226884 386092 226948
rect 386156 226884 386157 226948
rect 386091 226883 386157 226884
rect 383515 222868 383581 222869
rect 383515 222804 383516 222868
rect 383580 222804 383581 222868
rect 383515 222803 383581 222804
rect 388486 218653 388546 239670
rect 391062 224365 391122 239670
rect 391059 224364 391125 224365
rect 391059 224300 391060 224364
rect 391124 224300 391125 224364
rect 391059 224299 391125 224300
rect 388483 218652 388549 218653
rect 388483 218588 388484 218652
rect 388548 218588 388549 218652
rect 388483 218587 388549 218588
rect 381123 215932 381189 215933
rect 381123 215868 381124 215932
rect 381188 215868 381189 215932
rect 381123 215867 381189 215868
rect 356651 214708 356717 214709
rect 356651 214644 356652 214708
rect 356716 214644 356717 214708
rect 356651 214643 356717 214644
rect 393638 214573 393698 239670
rect 395846 239670 395996 239730
rect 398384 239730 398444 240040
rect 400968 239730 401028 240040
rect 403416 239730 403476 240040
rect 405864 239730 405924 240040
rect 408448 239730 408508 240040
rect 425750 240010 425916 240040
rect 425856 239869 425916 240010
rect 441662 240005 441722 253539
rect 441659 240004 441725 240005
rect 441659 239940 441660 240004
rect 441724 239940 441725 240004
rect 441659 239939 441725 239940
rect 425853 239868 425919 239869
rect 425853 239804 425854 239868
rect 425918 239804 425919 239868
rect 425853 239803 425919 239804
rect 425856 239730 425916 239803
rect 398384 239670 398482 239730
rect 400968 239670 401058 239730
rect 403416 239670 403634 239730
rect 395846 228309 395906 239670
rect 395843 228308 395909 228309
rect 395843 228244 395844 228308
rect 395908 228244 395909 228308
rect 395843 228243 395909 228244
rect 398422 224229 398482 239670
rect 400998 232525 401058 239670
rect 400995 232524 401061 232525
rect 400995 232460 400996 232524
rect 401060 232460 401061 232524
rect 400995 232459 401061 232460
rect 398419 224228 398485 224229
rect 398419 224164 398420 224228
rect 398484 224164 398485 224228
rect 398419 224163 398485 224164
rect 403574 221509 403634 239670
rect 405782 239670 405924 239730
rect 408358 239670 408508 239730
rect 425838 239670 425916 239730
rect 405782 234290 405842 239670
rect 408358 236605 408418 239670
rect 425838 237965 425898 239670
rect 425835 237964 425901 237965
rect 425835 237900 425836 237964
rect 425900 237900 425901 237964
rect 425835 237899 425901 237900
rect 408355 236604 408421 236605
rect 408355 236540 408356 236604
rect 408420 236540 408421 236604
rect 408355 236539 408421 236540
rect 405598 234230 405842 234290
rect 405598 229805 405658 234230
rect 405595 229804 405661 229805
rect 405595 229740 405596 229804
rect 405660 229740 405661 229804
rect 405595 229739 405661 229740
rect 409761 228174 410081 228206
rect 409761 227938 409803 228174
rect 410039 227938 410081 228174
rect 409761 227854 410081 227938
rect 409761 227618 409803 227854
rect 410039 227618 410081 227854
rect 409761 227586 410081 227618
rect 417603 228174 417923 228206
rect 417603 227938 417645 228174
rect 417881 227938 417923 228174
rect 417603 227854 417923 227938
rect 417603 227618 417645 227854
rect 417881 227618 417923 227854
rect 417603 227586 417923 227618
rect 425445 228174 425765 228206
rect 425445 227938 425487 228174
rect 425723 227938 425765 228174
rect 425445 227854 425765 227938
rect 425445 227618 425487 227854
rect 425723 227618 425765 227854
rect 425445 227586 425765 227618
rect 433287 228174 433607 228206
rect 433287 227938 433329 228174
rect 433565 227938 433607 228174
rect 433287 227854 433607 227938
rect 433287 227618 433329 227854
rect 433565 227618 433607 227854
rect 433287 227586 433607 227618
rect 405840 224454 406160 224486
rect 405840 224218 405882 224454
rect 406118 224218 406160 224454
rect 405840 224134 406160 224218
rect 405840 223898 405882 224134
rect 406118 223898 406160 224134
rect 405840 223866 406160 223898
rect 413682 224454 414002 224486
rect 413682 224218 413724 224454
rect 413960 224218 414002 224454
rect 413682 224134 414002 224218
rect 413682 223898 413724 224134
rect 413960 223898 414002 224134
rect 413682 223866 414002 223898
rect 421524 224454 421844 224486
rect 421524 224218 421566 224454
rect 421802 224218 421844 224454
rect 421524 224134 421844 224218
rect 421524 223898 421566 224134
rect 421802 223898 421844 224134
rect 421524 223866 421844 223898
rect 429366 224454 429686 224486
rect 429366 224218 429408 224454
rect 429644 224218 429686 224454
rect 429366 224134 429686 224218
rect 429366 223898 429408 224134
rect 429644 223898 429686 224134
rect 429366 223866 429686 223898
rect 403571 221508 403637 221509
rect 403571 221444 403572 221508
rect 403636 221444 403637 221508
rect 403571 221443 403637 221444
rect 409761 218174 410081 218206
rect 409761 217938 409803 218174
rect 410039 217938 410081 218174
rect 409761 217854 410081 217938
rect 409761 217618 409803 217854
rect 410039 217618 410081 217854
rect 409761 217586 410081 217618
rect 417603 218174 417923 218206
rect 417603 217938 417645 218174
rect 417881 217938 417923 218174
rect 417603 217854 417923 217938
rect 417603 217618 417645 217854
rect 417881 217618 417923 217854
rect 417603 217586 417923 217618
rect 425445 218174 425765 218206
rect 425445 217938 425487 218174
rect 425723 217938 425765 218174
rect 425445 217854 425765 217938
rect 425445 217618 425487 217854
rect 425723 217618 425765 217854
rect 425445 217586 425765 217618
rect 433287 218174 433607 218206
rect 433287 217938 433329 218174
rect 433565 217938 433607 218174
rect 433287 217854 433607 217938
rect 433287 217618 433329 217854
rect 433565 217618 433607 217854
rect 433287 217586 433607 217618
rect 393635 214572 393701 214573
rect 393635 214508 393636 214572
rect 393700 214508 393701 214572
rect 393635 214507 393701 214508
rect 405840 214454 406160 214486
rect 405840 214218 405882 214454
rect 406118 214218 406160 214454
rect 405840 214134 406160 214218
rect 405840 213898 405882 214134
rect 406118 213898 406160 214134
rect 405840 213866 406160 213898
rect 413682 214454 414002 214486
rect 413682 214218 413724 214454
rect 413960 214218 414002 214454
rect 413682 214134 414002 214218
rect 413682 213898 413724 214134
rect 413960 213898 414002 214134
rect 413682 213866 414002 213898
rect 421524 214454 421844 214486
rect 421524 214218 421566 214454
rect 421802 214218 421844 214454
rect 421524 214134 421844 214218
rect 421524 213898 421566 214134
rect 421802 213898 421844 214134
rect 421524 213866 421844 213898
rect 429366 214454 429686 214486
rect 429366 214218 429408 214454
rect 429644 214218 429686 214454
rect 429366 214134 429686 214218
rect 429366 213898 429408 214134
rect 429644 213898 429686 214134
rect 429366 213866 429686 213898
rect 341497 208174 341817 208206
rect 341497 207938 341539 208174
rect 341775 207938 341817 208174
rect 341497 207854 341817 207938
rect 341497 207618 341539 207854
rect 341775 207618 341817 207854
rect 341497 207586 341817 207618
rect 349339 208174 349659 208206
rect 349339 207938 349381 208174
rect 349617 207938 349659 208174
rect 349339 207854 349659 207938
rect 349339 207618 349381 207854
rect 349617 207618 349659 207854
rect 349339 207586 349659 207618
rect 357181 208174 357501 208206
rect 357181 207938 357223 208174
rect 357459 207938 357501 208174
rect 357181 207854 357501 207938
rect 357181 207618 357223 207854
rect 357459 207618 357501 207854
rect 357181 207586 357501 207618
rect 365023 208174 365343 208206
rect 365023 207938 365065 208174
rect 365301 207938 365343 208174
rect 365023 207854 365343 207938
rect 365023 207618 365065 207854
rect 365301 207618 365343 207854
rect 365023 207586 365343 207618
rect 375629 208174 375949 208206
rect 375629 207938 375671 208174
rect 375907 207938 375949 208174
rect 375629 207854 375949 207938
rect 375629 207618 375671 207854
rect 375907 207618 375949 207854
rect 375629 207586 375949 207618
rect 383471 208174 383791 208206
rect 383471 207938 383513 208174
rect 383749 207938 383791 208174
rect 383471 207854 383791 207938
rect 383471 207618 383513 207854
rect 383749 207618 383791 207854
rect 383471 207586 383791 207618
rect 391313 208174 391633 208206
rect 391313 207938 391355 208174
rect 391591 207938 391633 208174
rect 391313 207854 391633 207938
rect 391313 207618 391355 207854
rect 391591 207618 391633 207854
rect 391313 207586 391633 207618
rect 399155 208174 399475 208206
rect 399155 207938 399197 208174
rect 399433 207938 399475 208174
rect 399155 207854 399475 207938
rect 399155 207618 399197 207854
rect 399433 207618 399475 207854
rect 399155 207586 399475 207618
rect 409761 208174 410081 208206
rect 409761 207938 409803 208174
rect 410039 207938 410081 208174
rect 409761 207854 410081 207938
rect 409761 207618 409803 207854
rect 410039 207618 410081 207854
rect 409761 207586 410081 207618
rect 417603 208174 417923 208206
rect 417603 207938 417645 208174
rect 417881 207938 417923 208174
rect 417603 207854 417923 207938
rect 417603 207618 417645 207854
rect 417881 207618 417923 207854
rect 417603 207586 417923 207618
rect 425445 208174 425765 208206
rect 425445 207938 425487 208174
rect 425723 207938 425765 208174
rect 425445 207854 425765 207938
rect 425445 207618 425487 207854
rect 425723 207618 425765 207854
rect 425445 207586 425765 207618
rect 433287 208174 433607 208206
rect 433287 207938 433329 208174
rect 433565 207938 433607 208174
rect 433287 207854 433607 207938
rect 433287 207618 433329 207854
rect 433565 207618 433607 207854
rect 433287 207586 433607 207618
rect 443893 208174 444213 208206
rect 443893 207938 443935 208174
rect 444171 207938 444213 208174
rect 443893 207854 444213 207938
rect 443893 207618 443935 207854
rect 444171 207618 444213 207854
rect 443893 207586 444213 207618
rect 451735 208174 452055 208206
rect 451735 207938 451777 208174
rect 452013 207938 452055 208174
rect 451735 207854 452055 207938
rect 451735 207618 451777 207854
rect 452013 207618 452055 207854
rect 451735 207586 452055 207618
rect 459577 208174 459897 208206
rect 459577 207938 459619 208174
rect 459855 207938 459897 208174
rect 459577 207854 459897 207938
rect 459577 207618 459619 207854
rect 459855 207618 459897 207854
rect 459577 207586 459897 207618
rect 467419 208174 467739 208206
rect 467419 207938 467461 208174
rect 467697 207938 467739 208174
rect 467419 207854 467739 207938
rect 467419 207618 467461 207854
rect 467697 207618 467739 207854
rect 467419 207586 467739 207618
rect 478025 208174 478345 208206
rect 478025 207938 478067 208174
rect 478303 207938 478345 208174
rect 478025 207854 478345 207938
rect 478025 207618 478067 207854
rect 478303 207618 478345 207854
rect 478025 207586 478345 207618
rect 485867 208174 486187 208206
rect 485867 207938 485909 208174
rect 486145 207938 486187 208174
rect 485867 207854 486187 207938
rect 485867 207618 485909 207854
rect 486145 207618 486187 207854
rect 485867 207586 486187 207618
rect 493709 208174 494029 208206
rect 493709 207938 493751 208174
rect 493987 207938 494029 208174
rect 493709 207854 494029 207938
rect 493709 207618 493751 207854
rect 493987 207618 494029 207854
rect 493709 207586 494029 207618
rect 501551 208174 501871 208206
rect 501551 207938 501593 208174
rect 501829 207938 501871 208174
rect 501551 207854 501871 207938
rect 501551 207618 501593 207854
rect 501829 207618 501871 207854
rect 501551 207586 501871 207618
rect 512157 208174 512477 208206
rect 512157 207938 512199 208174
rect 512435 207938 512477 208174
rect 512157 207854 512477 207938
rect 512157 207618 512199 207854
rect 512435 207618 512477 207854
rect 512157 207586 512477 207618
rect 519999 208174 520319 208206
rect 519999 207938 520041 208174
rect 520277 207938 520319 208174
rect 519999 207854 520319 207938
rect 519999 207618 520041 207854
rect 520277 207618 520319 207854
rect 519999 207586 520319 207618
rect 527841 208174 528161 208206
rect 527841 207938 527883 208174
rect 528119 207938 528161 208174
rect 527841 207854 528161 207938
rect 527841 207618 527883 207854
rect 528119 207618 528161 207854
rect 527841 207586 528161 207618
rect 535683 208174 536003 208206
rect 535683 207938 535725 208174
rect 535961 207938 536003 208174
rect 535683 207854 536003 207938
rect 535683 207618 535725 207854
rect 535961 207618 536003 207854
rect 535683 207586 536003 207618
rect 546289 208174 546609 208206
rect 546289 207938 546331 208174
rect 546567 207938 546609 208174
rect 546289 207854 546609 207938
rect 546289 207618 546331 207854
rect 546567 207618 546609 207854
rect 546289 207586 546609 207618
rect 554131 208174 554451 208206
rect 554131 207938 554173 208174
rect 554409 207938 554451 208174
rect 554131 207854 554451 207938
rect 554131 207618 554173 207854
rect 554409 207618 554451 207854
rect 554131 207586 554451 207618
rect 561973 208174 562293 208206
rect 561973 207938 562015 208174
rect 562251 207938 562293 208174
rect 561973 207854 562293 207938
rect 561973 207618 562015 207854
rect 562251 207618 562293 207854
rect 561973 207586 562293 207618
rect 569815 208174 570135 208206
rect 569815 207938 569857 208174
rect 570093 207938 570135 208174
rect 569815 207854 570135 207938
rect 569815 207618 569857 207854
rect 570093 207618 570135 207854
rect 569815 207586 570135 207618
rect 337576 204454 337896 204486
rect 337576 204218 337618 204454
rect 337854 204218 337896 204454
rect 337576 204134 337896 204218
rect 337576 203898 337618 204134
rect 337854 203898 337896 204134
rect 337576 203866 337896 203898
rect 345418 204454 345738 204486
rect 345418 204218 345460 204454
rect 345696 204218 345738 204454
rect 345418 204134 345738 204218
rect 345418 203898 345460 204134
rect 345696 203898 345738 204134
rect 345418 203866 345738 203898
rect 353260 204454 353580 204486
rect 353260 204218 353302 204454
rect 353538 204218 353580 204454
rect 353260 204134 353580 204218
rect 353260 203898 353302 204134
rect 353538 203898 353580 204134
rect 353260 203866 353580 203898
rect 361102 204454 361422 204486
rect 361102 204218 361144 204454
rect 361380 204218 361422 204454
rect 361102 204134 361422 204218
rect 361102 203898 361144 204134
rect 361380 203898 361422 204134
rect 361102 203866 361422 203898
rect 371708 204454 372028 204486
rect 371708 204218 371750 204454
rect 371986 204218 372028 204454
rect 371708 204134 372028 204218
rect 371708 203898 371750 204134
rect 371986 203898 372028 204134
rect 371708 203866 372028 203898
rect 379550 204454 379870 204486
rect 379550 204218 379592 204454
rect 379828 204218 379870 204454
rect 379550 204134 379870 204218
rect 379550 203898 379592 204134
rect 379828 203898 379870 204134
rect 379550 203866 379870 203898
rect 387392 204454 387712 204486
rect 387392 204218 387434 204454
rect 387670 204218 387712 204454
rect 387392 204134 387712 204218
rect 387392 203898 387434 204134
rect 387670 203898 387712 204134
rect 387392 203866 387712 203898
rect 395234 204454 395554 204486
rect 395234 204218 395276 204454
rect 395512 204218 395554 204454
rect 395234 204134 395554 204218
rect 395234 203898 395276 204134
rect 395512 203898 395554 204134
rect 395234 203866 395554 203898
rect 405840 204454 406160 204486
rect 405840 204218 405882 204454
rect 406118 204218 406160 204454
rect 405840 204134 406160 204218
rect 405840 203898 405882 204134
rect 406118 203898 406160 204134
rect 405840 203866 406160 203898
rect 413682 204454 414002 204486
rect 413682 204218 413724 204454
rect 413960 204218 414002 204454
rect 413682 204134 414002 204218
rect 413682 203898 413724 204134
rect 413960 203898 414002 204134
rect 413682 203866 414002 203898
rect 421524 204454 421844 204486
rect 421524 204218 421566 204454
rect 421802 204218 421844 204454
rect 421524 204134 421844 204218
rect 421524 203898 421566 204134
rect 421802 203898 421844 204134
rect 421524 203866 421844 203898
rect 429366 204454 429686 204486
rect 429366 204218 429408 204454
rect 429644 204218 429686 204454
rect 429366 204134 429686 204218
rect 429366 203898 429408 204134
rect 429644 203898 429686 204134
rect 429366 203866 429686 203898
rect 439972 204454 440292 204486
rect 439972 204218 440014 204454
rect 440250 204218 440292 204454
rect 439972 204134 440292 204218
rect 439972 203898 440014 204134
rect 440250 203898 440292 204134
rect 439972 203866 440292 203898
rect 447814 204454 448134 204486
rect 447814 204218 447856 204454
rect 448092 204218 448134 204454
rect 447814 204134 448134 204218
rect 447814 203898 447856 204134
rect 448092 203898 448134 204134
rect 447814 203866 448134 203898
rect 455656 204454 455976 204486
rect 455656 204218 455698 204454
rect 455934 204218 455976 204454
rect 455656 204134 455976 204218
rect 455656 203898 455698 204134
rect 455934 203898 455976 204134
rect 455656 203866 455976 203898
rect 463498 204454 463818 204486
rect 463498 204218 463540 204454
rect 463776 204218 463818 204454
rect 463498 204134 463818 204218
rect 463498 203898 463540 204134
rect 463776 203898 463818 204134
rect 463498 203866 463818 203898
rect 474104 204454 474424 204486
rect 474104 204218 474146 204454
rect 474382 204218 474424 204454
rect 474104 204134 474424 204218
rect 474104 203898 474146 204134
rect 474382 203898 474424 204134
rect 474104 203866 474424 203898
rect 481946 204454 482266 204486
rect 481946 204218 481988 204454
rect 482224 204218 482266 204454
rect 481946 204134 482266 204218
rect 481946 203898 481988 204134
rect 482224 203898 482266 204134
rect 481946 203866 482266 203898
rect 489788 204454 490108 204486
rect 489788 204218 489830 204454
rect 490066 204218 490108 204454
rect 489788 204134 490108 204218
rect 489788 203898 489830 204134
rect 490066 203898 490108 204134
rect 489788 203866 490108 203898
rect 497630 204454 497950 204486
rect 497630 204218 497672 204454
rect 497908 204218 497950 204454
rect 497630 204134 497950 204218
rect 497630 203898 497672 204134
rect 497908 203898 497950 204134
rect 497630 203866 497950 203898
rect 508236 204454 508556 204486
rect 508236 204218 508278 204454
rect 508514 204218 508556 204454
rect 508236 204134 508556 204218
rect 508236 203898 508278 204134
rect 508514 203898 508556 204134
rect 508236 203866 508556 203898
rect 516078 204454 516398 204486
rect 516078 204218 516120 204454
rect 516356 204218 516398 204454
rect 516078 204134 516398 204218
rect 516078 203898 516120 204134
rect 516356 203898 516398 204134
rect 516078 203866 516398 203898
rect 523920 204454 524240 204486
rect 523920 204218 523962 204454
rect 524198 204218 524240 204454
rect 523920 204134 524240 204218
rect 523920 203898 523962 204134
rect 524198 203898 524240 204134
rect 523920 203866 524240 203898
rect 531762 204454 532082 204486
rect 531762 204218 531804 204454
rect 532040 204218 532082 204454
rect 531762 204134 532082 204218
rect 531762 203898 531804 204134
rect 532040 203898 532082 204134
rect 531762 203866 532082 203898
rect 542368 204454 542688 204486
rect 542368 204218 542410 204454
rect 542646 204218 542688 204454
rect 542368 204134 542688 204218
rect 542368 203898 542410 204134
rect 542646 203898 542688 204134
rect 542368 203866 542688 203898
rect 550210 204454 550530 204486
rect 550210 204218 550252 204454
rect 550488 204218 550530 204454
rect 550210 204134 550530 204218
rect 550210 203898 550252 204134
rect 550488 203898 550530 204134
rect 550210 203866 550530 203898
rect 558052 204454 558372 204486
rect 558052 204218 558094 204454
rect 558330 204218 558372 204454
rect 558052 204134 558372 204218
rect 558052 203898 558094 204134
rect 558330 203898 558372 204134
rect 558052 203866 558372 203898
rect 565894 204454 566214 204486
rect 565894 204218 565936 204454
rect 566172 204218 566214 204454
rect 565894 204134 566214 204218
rect 565894 203898 565936 204134
rect 566172 203898 566214 204134
rect 565894 203866 566214 203898
rect 341497 198174 341817 198206
rect 341497 197938 341539 198174
rect 341775 197938 341817 198174
rect 341497 197854 341817 197938
rect 341497 197618 341539 197854
rect 341775 197618 341817 197854
rect 341497 197586 341817 197618
rect 349339 198174 349659 198206
rect 349339 197938 349381 198174
rect 349617 197938 349659 198174
rect 349339 197854 349659 197938
rect 349339 197618 349381 197854
rect 349617 197618 349659 197854
rect 349339 197586 349659 197618
rect 357181 198174 357501 198206
rect 357181 197938 357223 198174
rect 357459 197938 357501 198174
rect 357181 197854 357501 197938
rect 357181 197618 357223 197854
rect 357459 197618 357501 197854
rect 357181 197586 357501 197618
rect 365023 198174 365343 198206
rect 365023 197938 365065 198174
rect 365301 197938 365343 198174
rect 365023 197854 365343 197938
rect 365023 197618 365065 197854
rect 365301 197618 365343 197854
rect 365023 197586 365343 197618
rect 375629 198174 375949 198206
rect 375629 197938 375671 198174
rect 375907 197938 375949 198174
rect 375629 197854 375949 197938
rect 375629 197618 375671 197854
rect 375907 197618 375949 197854
rect 375629 197586 375949 197618
rect 383471 198174 383791 198206
rect 383471 197938 383513 198174
rect 383749 197938 383791 198174
rect 383471 197854 383791 197938
rect 383471 197618 383513 197854
rect 383749 197618 383791 197854
rect 383471 197586 383791 197618
rect 391313 198174 391633 198206
rect 391313 197938 391355 198174
rect 391591 197938 391633 198174
rect 391313 197854 391633 197938
rect 391313 197618 391355 197854
rect 391591 197618 391633 197854
rect 391313 197586 391633 197618
rect 399155 198174 399475 198206
rect 399155 197938 399197 198174
rect 399433 197938 399475 198174
rect 399155 197854 399475 197938
rect 399155 197618 399197 197854
rect 399433 197618 399475 197854
rect 399155 197586 399475 197618
rect 409761 198174 410081 198206
rect 409761 197938 409803 198174
rect 410039 197938 410081 198174
rect 409761 197854 410081 197938
rect 409761 197618 409803 197854
rect 410039 197618 410081 197854
rect 409761 197586 410081 197618
rect 417603 198174 417923 198206
rect 417603 197938 417645 198174
rect 417881 197938 417923 198174
rect 417603 197854 417923 197938
rect 417603 197618 417645 197854
rect 417881 197618 417923 197854
rect 417603 197586 417923 197618
rect 425445 198174 425765 198206
rect 425445 197938 425487 198174
rect 425723 197938 425765 198174
rect 425445 197854 425765 197938
rect 425445 197618 425487 197854
rect 425723 197618 425765 197854
rect 425445 197586 425765 197618
rect 433287 198174 433607 198206
rect 433287 197938 433329 198174
rect 433565 197938 433607 198174
rect 433287 197854 433607 197938
rect 433287 197618 433329 197854
rect 433565 197618 433607 197854
rect 433287 197586 433607 197618
rect 443893 198174 444213 198206
rect 443893 197938 443935 198174
rect 444171 197938 444213 198174
rect 443893 197854 444213 197938
rect 443893 197618 443935 197854
rect 444171 197618 444213 197854
rect 443893 197586 444213 197618
rect 451735 198174 452055 198206
rect 451735 197938 451777 198174
rect 452013 197938 452055 198174
rect 451735 197854 452055 197938
rect 451735 197618 451777 197854
rect 452013 197618 452055 197854
rect 451735 197586 452055 197618
rect 459577 198174 459897 198206
rect 459577 197938 459619 198174
rect 459855 197938 459897 198174
rect 459577 197854 459897 197938
rect 459577 197618 459619 197854
rect 459855 197618 459897 197854
rect 459577 197586 459897 197618
rect 467419 198174 467739 198206
rect 467419 197938 467461 198174
rect 467697 197938 467739 198174
rect 467419 197854 467739 197938
rect 467419 197618 467461 197854
rect 467697 197618 467739 197854
rect 467419 197586 467739 197618
rect 478025 198174 478345 198206
rect 478025 197938 478067 198174
rect 478303 197938 478345 198174
rect 478025 197854 478345 197938
rect 478025 197618 478067 197854
rect 478303 197618 478345 197854
rect 478025 197586 478345 197618
rect 485867 198174 486187 198206
rect 485867 197938 485909 198174
rect 486145 197938 486187 198174
rect 485867 197854 486187 197938
rect 485867 197618 485909 197854
rect 486145 197618 486187 197854
rect 485867 197586 486187 197618
rect 493709 198174 494029 198206
rect 493709 197938 493751 198174
rect 493987 197938 494029 198174
rect 493709 197854 494029 197938
rect 493709 197618 493751 197854
rect 493987 197618 494029 197854
rect 493709 197586 494029 197618
rect 501551 198174 501871 198206
rect 501551 197938 501593 198174
rect 501829 197938 501871 198174
rect 501551 197854 501871 197938
rect 501551 197618 501593 197854
rect 501829 197618 501871 197854
rect 501551 197586 501871 197618
rect 512157 198174 512477 198206
rect 512157 197938 512199 198174
rect 512435 197938 512477 198174
rect 512157 197854 512477 197938
rect 512157 197618 512199 197854
rect 512435 197618 512477 197854
rect 512157 197586 512477 197618
rect 519999 198174 520319 198206
rect 519999 197938 520041 198174
rect 520277 197938 520319 198174
rect 519999 197854 520319 197938
rect 519999 197618 520041 197854
rect 520277 197618 520319 197854
rect 519999 197586 520319 197618
rect 527841 198174 528161 198206
rect 527841 197938 527883 198174
rect 528119 197938 528161 198174
rect 527841 197854 528161 197938
rect 527841 197618 527883 197854
rect 528119 197618 528161 197854
rect 527841 197586 528161 197618
rect 535683 198174 536003 198206
rect 535683 197938 535725 198174
rect 535961 197938 536003 198174
rect 535683 197854 536003 197938
rect 535683 197618 535725 197854
rect 535961 197618 536003 197854
rect 535683 197586 536003 197618
rect 546289 198174 546609 198206
rect 546289 197938 546331 198174
rect 546567 197938 546609 198174
rect 546289 197854 546609 197938
rect 546289 197618 546331 197854
rect 546567 197618 546609 197854
rect 546289 197586 546609 197618
rect 554131 198174 554451 198206
rect 554131 197938 554173 198174
rect 554409 197938 554451 198174
rect 554131 197854 554451 197938
rect 554131 197618 554173 197854
rect 554409 197618 554451 197854
rect 554131 197586 554451 197618
rect 561973 198174 562293 198206
rect 561973 197938 562015 198174
rect 562251 197938 562293 198174
rect 561973 197854 562293 197938
rect 561973 197618 562015 197854
rect 562251 197618 562293 197854
rect 561973 197586 562293 197618
rect 569815 198174 570135 198206
rect 569815 197938 569857 198174
rect 570093 197938 570135 198174
rect 569815 197854 570135 197938
rect 569815 197618 569857 197854
rect 570093 197618 570135 197854
rect 569815 197586 570135 197618
rect 337576 194454 337896 194486
rect 337576 194218 337618 194454
rect 337854 194218 337896 194454
rect 337576 194134 337896 194218
rect 337576 193898 337618 194134
rect 337854 193898 337896 194134
rect 337576 193866 337896 193898
rect 345418 194454 345738 194486
rect 345418 194218 345460 194454
rect 345696 194218 345738 194454
rect 345418 194134 345738 194218
rect 345418 193898 345460 194134
rect 345696 193898 345738 194134
rect 345418 193866 345738 193898
rect 353260 194454 353580 194486
rect 353260 194218 353302 194454
rect 353538 194218 353580 194454
rect 353260 194134 353580 194218
rect 353260 193898 353302 194134
rect 353538 193898 353580 194134
rect 353260 193866 353580 193898
rect 361102 194454 361422 194486
rect 361102 194218 361144 194454
rect 361380 194218 361422 194454
rect 361102 194134 361422 194218
rect 361102 193898 361144 194134
rect 361380 193898 361422 194134
rect 361102 193866 361422 193898
rect 371708 194454 372028 194486
rect 371708 194218 371750 194454
rect 371986 194218 372028 194454
rect 371708 194134 372028 194218
rect 371708 193898 371750 194134
rect 371986 193898 372028 194134
rect 371708 193866 372028 193898
rect 379550 194454 379870 194486
rect 379550 194218 379592 194454
rect 379828 194218 379870 194454
rect 379550 194134 379870 194218
rect 379550 193898 379592 194134
rect 379828 193898 379870 194134
rect 379550 193866 379870 193898
rect 387392 194454 387712 194486
rect 387392 194218 387434 194454
rect 387670 194218 387712 194454
rect 387392 194134 387712 194218
rect 387392 193898 387434 194134
rect 387670 193898 387712 194134
rect 387392 193866 387712 193898
rect 395234 194454 395554 194486
rect 395234 194218 395276 194454
rect 395512 194218 395554 194454
rect 395234 194134 395554 194218
rect 395234 193898 395276 194134
rect 395512 193898 395554 194134
rect 395234 193866 395554 193898
rect 405840 194454 406160 194486
rect 405840 194218 405882 194454
rect 406118 194218 406160 194454
rect 405840 194134 406160 194218
rect 405840 193898 405882 194134
rect 406118 193898 406160 194134
rect 405840 193866 406160 193898
rect 413682 194454 414002 194486
rect 413682 194218 413724 194454
rect 413960 194218 414002 194454
rect 413682 194134 414002 194218
rect 413682 193898 413724 194134
rect 413960 193898 414002 194134
rect 413682 193866 414002 193898
rect 421524 194454 421844 194486
rect 421524 194218 421566 194454
rect 421802 194218 421844 194454
rect 421524 194134 421844 194218
rect 421524 193898 421566 194134
rect 421802 193898 421844 194134
rect 421524 193866 421844 193898
rect 429366 194454 429686 194486
rect 429366 194218 429408 194454
rect 429644 194218 429686 194454
rect 429366 194134 429686 194218
rect 429366 193898 429408 194134
rect 429644 193898 429686 194134
rect 429366 193866 429686 193898
rect 439972 194454 440292 194486
rect 439972 194218 440014 194454
rect 440250 194218 440292 194454
rect 439972 194134 440292 194218
rect 439972 193898 440014 194134
rect 440250 193898 440292 194134
rect 439972 193866 440292 193898
rect 447814 194454 448134 194486
rect 447814 194218 447856 194454
rect 448092 194218 448134 194454
rect 447814 194134 448134 194218
rect 447814 193898 447856 194134
rect 448092 193898 448134 194134
rect 447814 193866 448134 193898
rect 455656 194454 455976 194486
rect 455656 194218 455698 194454
rect 455934 194218 455976 194454
rect 455656 194134 455976 194218
rect 455656 193898 455698 194134
rect 455934 193898 455976 194134
rect 455656 193866 455976 193898
rect 463498 194454 463818 194486
rect 463498 194218 463540 194454
rect 463776 194218 463818 194454
rect 463498 194134 463818 194218
rect 463498 193898 463540 194134
rect 463776 193898 463818 194134
rect 463498 193866 463818 193898
rect 474104 194454 474424 194486
rect 474104 194218 474146 194454
rect 474382 194218 474424 194454
rect 474104 194134 474424 194218
rect 474104 193898 474146 194134
rect 474382 193898 474424 194134
rect 474104 193866 474424 193898
rect 481946 194454 482266 194486
rect 481946 194218 481988 194454
rect 482224 194218 482266 194454
rect 481946 194134 482266 194218
rect 481946 193898 481988 194134
rect 482224 193898 482266 194134
rect 481946 193866 482266 193898
rect 489788 194454 490108 194486
rect 489788 194218 489830 194454
rect 490066 194218 490108 194454
rect 489788 194134 490108 194218
rect 489788 193898 489830 194134
rect 490066 193898 490108 194134
rect 489788 193866 490108 193898
rect 497630 194454 497950 194486
rect 497630 194218 497672 194454
rect 497908 194218 497950 194454
rect 497630 194134 497950 194218
rect 497630 193898 497672 194134
rect 497908 193898 497950 194134
rect 497630 193866 497950 193898
rect 508236 194454 508556 194486
rect 508236 194218 508278 194454
rect 508514 194218 508556 194454
rect 508236 194134 508556 194218
rect 508236 193898 508278 194134
rect 508514 193898 508556 194134
rect 508236 193866 508556 193898
rect 516078 194454 516398 194486
rect 516078 194218 516120 194454
rect 516356 194218 516398 194454
rect 516078 194134 516398 194218
rect 516078 193898 516120 194134
rect 516356 193898 516398 194134
rect 516078 193866 516398 193898
rect 523920 194454 524240 194486
rect 523920 194218 523962 194454
rect 524198 194218 524240 194454
rect 523920 194134 524240 194218
rect 523920 193898 523962 194134
rect 524198 193898 524240 194134
rect 523920 193866 524240 193898
rect 531762 194454 532082 194486
rect 531762 194218 531804 194454
rect 532040 194218 532082 194454
rect 531762 194134 532082 194218
rect 531762 193898 531804 194134
rect 532040 193898 532082 194134
rect 531762 193866 532082 193898
rect 542368 194454 542688 194486
rect 542368 194218 542410 194454
rect 542646 194218 542688 194454
rect 542368 194134 542688 194218
rect 542368 193898 542410 194134
rect 542646 193898 542688 194134
rect 542368 193866 542688 193898
rect 550210 194454 550530 194486
rect 550210 194218 550252 194454
rect 550488 194218 550530 194454
rect 550210 194134 550530 194218
rect 550210 193898 550252 194134
rect 550488 193898 550530 194134
rect 550210 193866 550530 193898
rect 558052 194454 558372 194486
rect 558052 194218 558094 194454
rect 558330 194218 558372 194454
rect 558052 194134 558372 194218
rect 558052 193898 558094 194134
rect 558330 193898 558372 194134
rect 558052 193866 558372 193898
rect 565894 194454 566214 194486
rect 565894 194218 565936 194454
rect 566172 194218 566214 194454
rect 565894 194134 566214 194218
rect 565894 193898 565936 194134
rect 566172 193898 566214 194134
rect 565894 193866 566214 193898
rect 301083 191860 301149 191861
rect 301083 191796 301084 191860
rect 301148 191796 301149 191860
rect 301083 191795 301149 191796
rect 335123 191860 335189 191861
rect 335123 191796 335124 191860
rect 335188 191796 335189 191860
rect 335123 191795 335189 191796
rect 337331 191860 337397 191861
rect 337331 191796 337332 191860
rect 337396 191796 337397 191860
rect 337331 191795 337397 191796
rect 298691 190772 298757 190773
rect 298691 190708 298692 190772
rect 298756 190708 298757 190772
rect 298691 190707 298757 190708
rect 298694 190501 298754 190707
rect 298691 190500 298757 190501
rect 298691 190436 298692 190500
rect 298756 190436 298757 190500
rect 298691 190435 298757 190436
rect 296851 188596 296917 188597
rect 296851 188532 296852 188596
rect 296916 188532 296917 188596
rect 296851 188531 296917 188532
rect 296854 186013 296914 188531
rect 297955 186828 298021 186829
rect 297955 186764 297956 186828
rect 298020 186764 298021 186828
rect 297955 186763 298021 186764
rect 297403 186692 297469 186693
rect 297403 186628 297404 186692
rect 297468 186628 297469 186692
rect 297403 186627 297469 186628
rect 296851 186012 296917 186013
rect 296851 185948 296852 186012
rect 296916 185948 296917 186012
rect 296851 185947 296917 185948
rect 296854 180437 296914 185947
rect 296851 180436 296917 180437
rect 296851 180372 296852 180436
rect 296916 180372 296917 180436
rect 296851 180371 296917 180372
rect 296667 176628 296733 176629
rect 296667 176564 296668 176628
rect 296732 176564 296733 176628
rect 296667 176563 296733 176564
rect 296670 167109 296730 176563
rect 296667 167108 296733 167109
rect 296667 167044 296668 167108
rect 296732 167044 296733 167108
rect 296667 167043 296733 167044
rect 296667 161532 296733 161533
rect 296667 161468 296668 161532
rect 296732 161468 296733 161532
rect 296667 161467 296733 161468
rect 296670 161261 296730 161467
rect 296667 161260 296733 161261
rect 296667 161196 296668 161260
rect 296732 161196 296733 161260
rect 296667 161195 296733 161196
rect 296483 156908 296549 156909
rect 296483 156844 296484 156908
rect 296548 156844 296549 156908
rect 296483 156843 296549 156844
rect 296667 151876 296733 151877
rect 296667 151830 296668 151876
rect 296486 151812 296668 151830
rect 296732 151812 296733 151876
rect 296486 151811 296733 151812
rect 296486 151770 296730 151811
rect 296486 66330 296546 151770
rect 297035 67556 297101 67557
rect 297035 67492 297036 67556
rect 297100 67492 297101 67556
rect 297035 67491 297101 67492
rect 296486 66270 296730 66330
rect 296670 65620 296730 66270
rect 297038 65620 297098 67491
rect 297406 65620 297466 186627
rect 297958 186421 298018 186763
rect 298139 186556 298205 186557
rect 298139 186492 298140 186556
rect 298204 186492 298205 186556
rect 298139 186491 298205 186492
rect 297955 186420 298021 186421
rect 297955 186356 297956 186420
rect 298020 186356 298021 186420
rect 297955 186355 298021 186356
rect 297958 180810 298018 186355
rect 297774 180750 298018 180810
rect 297774 65620 297834 180750
rect 298142 65620 298202 186491
rect 298323 177444 298389 177445
rect 298323 177380 298324 177444
rect 298388 177380 298389 177444
rect 298323 177379 298389 177380
rect 298326 67557 298386 177379
rect 298323 67556 298389 67557
rect 298323 67492 298324 67556
rect 298388 67492 298389 67556
rect 298323 67491 298389 67492
rect 298694 66333 298754 190435
rect 299795 189684 299861 189685
rect 299795 189620 299796 189684
rect 299860 189620 299861 189684
rect 299795 189619 299861 189620
rect 299243 187644 299309 187645
rect 299243 187580 299244 187644
rect 299308 187580 299309 187644
rect 299243 187579 299309 187580
rect 298875 179756 298941 179757
rect 298875 179692 298876 179756
rect 298940 179692 298941 179756
rect 298875 179691 298941 179692
rect 298878 178669 298938 179691
rect 299246 179621 299306 187579
rect 299798 187237 299858 189619
rect 299979 189412 300045 189413
rect 299979 189348 299980 189412
rect 300044 189348 300045 189412
rect 299979 189347 300045 189348
rect 299982 187509 300042 189347
rect 300899 188324 300965 188325
rect 300899 188260 300900 188324
rect 300964 188260 300965 188324
rect 300899 188259 300965 188260
rect 299979 187508 300045 187509
rect 299979 187444 299980 187508
rect 300044 187444 300045 187508
rect 299979 187443 300045 187444
rect 299795 187236 299861 187237
rect 299795 187172 299796 187236
rect 299860 187172 299861 187236
rect 299795 187171 299861 187172
rect 299427 186692 299493 186693
rect 299427 186628 299428 186692
rect 299492 186628 299493 186692
rect 299427 186627 299493 186628
rect 299430 186285 299490 186627
rect 299427 186284 299493 186285
rect 299427 186220 299428 186284
rect 299492 186220 299493 186284
rect 299427 186219 299493 186220
rect 299795 185876 299861 185877
rect 299795 185812 299796 185876
rect 299860 185812 299861 185876
rect 299795 185811 299861 185812
rect 299243 179620 299309 179621
rect 299243 179556 299244 179620
rect 299308 179556 299309 179620
rect 299243 179555 299309 179556
rect 299798 178941 299858 185811
rect 299982 184653 300042 187443
rect 300163 187236 300229 187237
rect 300163 187172 300164 187236
rect 300228 187172 300229 187236
rect 300163 187171 300229 187172
rect 299979 184652 300045 184653
rect 299979 184588 299980 184652
rect 300044 184588 300045 184652
rect 299979 184587 300045 184588
rect 300166 180810 300226 187171
rect 300715 187100 300781 187101
rect 300715 187036 300716 187100
rect 300780 187036 300781 187100
rect 300715 187035 300781 187036
rect 300531 183836 300597 183837
rect 300531 183772 300532 183836
rect 300596 183772 300597 183836
rect 300531 183771 300597 183772
rect 299982 180750 300226 180810
rect 299795 178940 299861 178941
rect 299795 178876 299796 178940
rect 299860 178876 299861 178940
rect 299795 178875 299861 178876
rect 298875 178668 298941 178669
rect 298875 178604 298876 178668
rect 298940 178604 298941 178668
rect 298875 178603 298941 178604
rect 299795 71092 299861 71093
rect 299795 71028 299796 71092
rect 299860 71028 299861 71092
rect 299795 71027 299861 71028
rect 299243 67692 299309 67693
rect 299243 67628 299244 67692
rect 299308 67628 299309 67692
rect 299243 67627 299309 67628
rect 298875 67556 298941 67557
rect 298875 67492 298876 67556
rect 298940 67492 298941 67556
rect 298875 67491 298941 67492
rect 298878 66469 298938 67491
rect 298875 66468 298941 66469
rect 298875 66404 298876 66468
rect 298940 66404 298941 66468
rect 298875 66403 298941 66404
rect 298691 66332 298757 66333
rect 298691 66268 298692 66332
rect 298756 66268 298757 66332
rect 298691 66267 298757 66268
rect 298694 65650 298754 66267
rect 298540 65590 298754 65650
rect 298878 65620 298938 66403
rect 299246 65620 299306 67627
rect 299798 67557 299858 71027
rect 299982 67965 300042 180750
rect 300534 180301 300594 183771
rect 300531 180300 300597 180301
rect 300531 180236 300532 180300
rect 300596 180236 300597 180300
rect 300531 180235 300597 180236
rect 300163 180164 300229 180165
rect 300163 180100 300164 180164
rect 300228 180100 300229 180164
rect 300163 180099 300229 180100
rect 300166 68917 300226 180099
rect 300718 157045 300778 187035
rect 300902 184653 300962 188259
rect 301086 187917 301146 191795
rect 303570 190400 303630 191044
rect 304306 190400 304366 191420
rect 305042 190400 305102 191080
rect 305778 190400 305838 191080
rect 306514 190400 306574 191080
rect 307250 190400 307310 191080
rect 307986 190400 308046 191080
rect 308722 190400 308782 191080
rect 309458 190400 309518 191080
rect 310194 190400 310254 191080
rect 310930 190400 310990 191080
rect 311666 190400 311726 191080
rect 312402 190400 312462 191080
rect 313138 190400 313198 191080
rect 313874 190400 313934 191080
rect 314610 190400 314670 191080
rect 315346 190400 315406 191080
rect 316082 190400 316142 191080
rect 316818 190400 316878 191080
rect 317554 190400 317614 191420
rect 318290 190400 318350 191420
rect 319026 190400 319086 191080
rect 319762 190400 319822 191420
rect 320498 190400 320558 191420
rect 321234 190400 321294 191420
rect 321970 190400 322030 191420
rect 322706 190400 322766 191420
rect 323442 190400 323502 191080
rect 324178 190400 324238 191080
rect 324914 190400 324974 191080
rect 325650 190400 325710 191080
rect 326386 190400 326446 191080
rect 327122 190400 327182 191080
rect 327858 190400 327918 191080
rect 328594 190400 328654 191080
rect 329330 190400 329390 191080
rect 330066 190400 330126 191080
rect 330802 190400 330862 191080
rect 331538 190400 331598 191080
rect 332274 190400 332334 191080
rect 333010 190400 333070 191080
rect 333746 190400 333806 191080
rect 334482 190400 334542 191080
rect 335126 190470 335186 191795
rect 335126 190410 335278 190470
rect 335218 190400 335278 190410
rect 337702 190060 337762 191044
rect 338438 190400 338498 191080
rect 339174 190400 339234 191080
rect 339910 190060 339970 191080
rect 340646 190060 340706 191044
rect 341382 190400 341442 191044
rect 342118 190060 342178 191044
rect 342854 190400 342914 191044
rect 343590 190060 343650 191044
rect 344326 190060 344386 191044
rect 345062 190400 345122 191044
rect 345798 190060 345858 191080
rect 346534 190400 346594 191080
rect 347270 190400 347330 191080
rect 348006 190060 348066 191080
rect 348742 190060 348802 191080
rect 349478 190060 349538 191080
rect 350214 190060 350274 191080
rect 350950 190400 351010 191080
rect 351686 190400 351746 191080
rect 352422 190400 352482 191080
rect 353158 190400 353218 191080
rect 353894 190400 353954 191080
rect 354630 190400 354690 191080
rect 355366 190400 355426 191080
rect 356102 190400 356162 191080
rect 356838 190400 356898 191080
rect 357574 190400 357634 191080
rect 358310 190400 358370 191080
rect 359046 190400 359106 191080
rect 359782 190400 359842 191080
rect 360518 190400 360578 191420
rect 361254 190400 361314 191080
rect 361990 190400 362050 191080
rect 362726 190400 362786 191080
rect 363462 190400 363522 191080
rect 364198 190400 364258 191080
rect 364934 190400 364994 191080
rect 365670 190400 365730 191080
rect 366406 190400 366466 191420
rect 367142 190400 367202 191080
rect 367878 190400 367938 191080
rect 368614 190400 368674 191420
rect 371834 190400 371894 191044
rect 372570 190400 372630 191080
rect 373306 190400 373366 191080
rect 374042 190400 374102 191044
rect 374778 190400 374838 191044
rect 375514 190400 375574 191080
rect 376250 190400 376310 191080
rect 376986 190400 377046 191080
rect 377722 190400 377782 191080
rect 378458 190400 378518 191044
rect 379194 190400 379254 191044
rect 379930 190400 379990 191044
rect 380666 190400 380726 191044
rect 381402 190400 381462 191044
rect 382138 190400 382198 191044
rect 382874 190400 382934 191044
rect 383610 190400 383670 191044
rect 384346 190400 384406 191044
rect 385082 190400 385142 191044
rect 385818 190400 385878 191080
rect 386554 190400 386614 191080
rect 387290 190400 387350 191080
rect 388026 190400 388086 191080
rect 388762 190400 388822 191080
rect 389498 190400 389558 191080
rect 390234 190400 390294 191080
rect 390970 190400 391030 191080
rect 391706 190400 391766 191420
rect 392442 190400 392502 191080
rect 393178 190400 393238 191080
rect 393914 190400 393974 191420
rect 394650 190400 394710 191080
rect 395386 190400 395446 191080
rect 396122 190400 396182 191080
rect 396858 190400 396918 191080
rect 397594 190400 397654 191080
rect 398330 190400 398390 191080
rect 399066 190400 399126 191080
rect 399802 190400 399862 191080
rect 400538 190400 400598 191080
rect 401274 190400 401334 191080
rect 402010 190400 402070 191080
rect 402746 190770 402806 191420
rect 402654 190710 402806 190770
rect 402654 190470 402714 190710
rect 402654 190410 402806 190470
rect 402746 190400 402806 190410
rect 405966 190400 406026 191044
rect 406702 190400 406762 191420
rect 407438 190400 407498 191080
rect 408174 190060 408234 191080
rect 408910 190060 408970 191080
rect 409646 190060 409706 191080
rect 410382 190060 410442 191080
rect 411118 190060 411178 191080
rect 411854 190060 411914 191080
rect 412590 190060 412650 191080
rect 413326 190060 413386 191080
rect 414062 190060 414122 191080
rect 414798 190060 414858 191080
rect 415534 190060 415594 191080
rect 416270 190060 416330 191080
rect 417006 190060 417066 191044
rect 417742 190060 417802 191044
rect 418478 190400 418538 191044
rect 419214 190060 419274 191044
rect 419950 190400 420010 191080
rect 420686 190400 420746 191080
rect 421422 190400 421482 191080
rect 422158 190400 422218 191080
rect 422894 190400 422954 191080
rect 423630 190400 423690 191080
rect 424366 190400 424426 191080
rect 425102 190400 425162 191420
rect 425838 190400 425898 191080
rect 426574 190400 426634 191080
rect 427310 190400 427370 191080
rect 428046 190400 428106 191080
rect 428782 190400 428842 191080
rect 429518 190400 429578 191080
rect 430254 190400 430314 191080
rect 430990 190400 431050 191420
rect 431726 190400 431786 191080
rect 432462 190400 432522 191080
rect 433198 190400 433258 191080
rect 433934 190400 433994 191080
rect 434670 190400 434730 191080
rect 435406 190400 435466 191080
rect 436142 190400 436202 191080
rect 436878 190400 436938 191080
rect 440098 190400 440158 191044
rect 440834 190400 440894 191044
rect 441570 190400 441630 191044
rect 442306 190400 442366 191080
rect 443042 190400 443102 191080
rect 443778 190400 443838 191080
rect 444514 190400 444574 191080
rect 445250 190400 445310 191080
rect 445986 190400 446046 191044
rect 446722 190400 446782 191044
rect 447458 190400 447518 191080
rect 448194 190400 448254 191044
rect 448930 190400 448990 191044
rect 449666 190400 449726 191044
rect 450402 190400 450462 191044
rect 451138 190400 451198 191044
rect 451874 190400 451934 191044
rect 452610 190400 452670 191044
rect 453346 190400 453406 191044
rect 454082 190400 454142 191080
rect 454818 190400 454878 191080
rect 455554 190400 455614 191080
rect 456290 190400 456350 191080
rect 457026 190400 457086 191080
rect 457762 190400 457822 191080
rect 458498 190400 458558 191080
rect 459234 190400 459294 191080
rect 459970 190400 460030 191080
rect 460706 190400 460766 191080
rect 461442 190400 461502 191080
rect 462178 190400 462238 191080
rect 462914 190400 462974 191080
rect 463650 190400 463710 191080
rect 464386 190400 464446 191080
rect 465122 190400 465182 191080
rect 465858 190400 465918 191080
rect 466594 190400 466654 191080
rect 467330 190400 467390 191080
rect 468066 190400 468126 191080
rect 468802 190400 468862 191080
rect 469538 190400 469598 191080
rect 470274 190400 470334 191080
rect 471010 190400 471070 191080
rect 474230 190400 474290 191044
rect 474966 190400 475026 191420
rect 475702 190060 475762 191044
rect 476438 190400 476498 191044
rect 477174 190060 477234 191044
rect 477910 190060 477970 191044
rect 478646 190400 478706 191044
rect 479382 190400 479442 191044
rect 480118 190060 480178 191044
rect 480854 190060 480914 191080
rect 481590 190400 481650 191080
rect 482326 190400 482386 191044
rect 483062 190400 483122 191044
rect 483798 190400 483858 191044
rect 484534 190060 484594 191044
rect 485270 190400 485330 191044
rect 486006 190060 486066 191044
rect 486742 190400 486802 191044
rect 487478 190060 487538 191044
rect 488214 190400 488274 191080
rect 488950 190400 489010 191080
rect 489686 190400 489746 191080
rect 490422 190400 490482 191080
rect 491158 190400 491218 191080
rect 491894 190400 491954 191080
rect 492630 190400 492690 191080
rect 493366 190400 493426 191080
rect 494102 190400 494162 191080
rect 494838 190400 494898 191080
rect 495574 190400 495634 191080
rect 496310 190400 496370 191080
rect 497046 190400 497106 191080
rect 497782 190400 497842 191080
rect 498518 190400 498578 191080
rect 499254 190400 499314 191080
rect 499990 190060 500050 191080
rect 500726 190400 500786 191080
rect 501462 190060 501522 191080
rect 502198 190400 502258 191080
rect 502934 190400 502994 191080
rect 503670 190400 503730 191080
rect 504406 190400 504466 191080
rect 505142 190400 505202 191080
rect 508362 190400 508422 191044
rect 509098 190400 509158 191080
rect 509834 190400 509894 191044
rect 510570 190400 510630 191044
rect 511306 190400 511366 191080
rect 512042 190400 512102 191044
rect 512778 190400 512838 191080
rect 513514 190400 513574 191080
rect 514250 190400 514310 191080
rect 514986 190400 515046 191080
rect 515722 190400 515782 191080
rect 516458 190400 516518 191044
rect 517194 190400 517254 191044
rect 517930 190400 517990 191044
rect 518666 190400 518726 191044
rect 519402 190400 519462 191044
rect 520138 190400 520198 191044
rect 520874 190400 520934 191044
rect 521610 190400 521670 191044
rect 522346 190400 522406 191080
rect 523082 190400 523142 191080
rect 523818 190400 523878 191080
rect 524554 190400 524614 191080
rect 525290 190400 525350 191080
rect 526026 190400 526086 191080
rect 526762 190400 526822 191080
rect 527498 190400 527558 191080
rect 528234 190400 528294 191080
rect 528970 190400 529030 191080
rect 529706 190400 529766 191080
rect 530442 190400 530502 191080
rect 531178 190400 531238 191080
rect 531914 190400 531974 191080
rect 532650 190400 532710 191080
rect 533386 190400 533446 191080
rect 534122 190400 534182 191080
rect 534858 190400 534918 191080
rect 535594 190400 535654 191080
rect 536330 190400 536390 191080
rect 537066 190400 537126 191080
rect 537802 190400 537862 191080
rect 538538 190400 538598 191080
rect 539274 190400 539334 191080
rect 542494 190400 542554 191044
rect 543230 190400 543290 191044
rect 543966 190060 544026 191044
rect 544702 190400 544762 191080
rect 545438 190400 545498 191044
rect 546174 190060 546234 191044
rect 546910 190060 546970 191044
rect 547646 190060 547706 191080
rect 548382 190400 548442 191080
rect 549118 190400 549178 191080
rect 549854 190060 549914 191080
rect 550590 190400 550650 191044
rect 551326 190060 551386 191044
rect 552062 190060 552122 191044
rect 552798 190060 552858 191044
rect 553534 190060 553594 191044
rect 554270 190060 554330 191044
rect 555006 190400 555066 191044
rect 555742 190060 555802 191044
rect 556478 190400 556538 191080
rect 557214 190400 557274 191080
rect 557950 190400 558010 191080
rect 558686 190400 558746 191080
rect 559422 190400 559482 191080
rect 560158 190400 560218 191080
rect 560894 190400 560954 191080
rect 561630 190400 561690 191080
rect 562366 190400 562426 191080
rect 563102 190400 563162 191080
rect 563838 190400 563898 191080
rect 564574 190400 564634 191080
rect 565310 190400 565370 191080
rect 566046 190400 566106 191080
rect 566782 190400 566842 191080
rect 567518 190400 567578 191080
rect 568254 190400 568314 191080
rect 568990 190400 569050 191080
rect 569726 190400 569786 191080
rect 570462 190400 570522 191080
rect 571198 190400 571258 191080
rect 571934 190400 571994 191080
rect 572670 190400 572730 191080
rect 573406 190400 573466 191080
rect 302739 189004 302805 189005
rect 302739 188940 302740 189004
rect 302804 188940 302805 189004
rect 302739 188939 302805 188940
rect 302742 188869 302802 188939
rect 302739 188868 302805 188869
rect 302739 188804 302740 188868
rect 302804 188804 302805 188868
rect 302739 188803 302805 188804
rect 301267 188732 301333 188733
rect 301267 188668 301268 188732
rect 301332 188668 301333 188732
rect 301267 188667 301333 188668
rect 301083 187916 301149 187917
rect 301083 187852 301084 187916
rect 301148 187852 301149 187916
rect 301083 187851 301149 187852
rect 300899 184652 300965 184653
rect 300899 184588 300900 184652
rect 300964 184588 300965 184652
rect 300899 184587 300965 184588
rect 301083 182612 301149 182613
rect 301083 182548 301084 182612
rect 301148 182548 301149 182612
rect 301083 182547 301149 182548
rect 300899 182476 300965 182477
rect 300899 182412 300900 182476
rect 300964 182412 300965 182476
rect 300899 182411 300965 182412
rect 300902 179757 300962 182411
rect 300899 179756 300965 179757
rect 300899 179692 300900 179756
rect 300964 179692 300965 179756
rect 300899 179691 300965 179692
rect 301086 179213 301146 182547
rect 301270 182205 301330 188667
rect 302742 188325 302802 188803
rect 302739 188324 302805 188325
rect 302739 188260 302740 188324
rect 302804 188260 302805 188324
rect 302739 188259 302805 188260
rect 302463 188188 302529 188189
rect 302463 188124 302464 188188
rect 302528 188124 302529 188188
rect 302463 188123 302529 188124
rect 337147 188174 337467 188206
rect 302466 188050 302526 188123
rect 302374 187990 302526 188050
rect 301451 187916 301517 187917
rect 301451 187852 301452 187916
rect 301516 187852 301517 187916
rect 301451 187851 301517 187852
rect 301267 182204 301333 182205
rect 301267 182140 301268 182204
rect 301332 182140 301333 182204
rect 301267 182139 301333 182140
rect 301083 179212 301149 179213
rect 301083 179148 301084 179212
rect 301148 179148 301149 179212
rect 301083 179147 301149 179148
rect 300715 157044 300781 157045
rect 300715 156980 300716 157044
rect 300780 156980 300781 157044
rect 300715 156979 300781 156980
rect 300715 156636 300781 156637
rect 300715 156572 300716 156636
rect 300780 156572 300781 156636
rect 300715 156571 300781 156572
rect 300718 155410 300778 156571
rect 300718 155350 300962 155410
rect 300902 153781 300962 155350
rect 300899 153780 300965 153781
rect 300899 153716 300900 153780
rect 300964 153716 300965 153780
rect 300899 153715 300965 153716
rect 301454 74550 301514 187851
rect 301635 184380 301701 184381
rect 301635 184316 301636 184380
rect 301700 184316 301701 184380
rect 301635 184315 301701 184316
rect 301638 179077 301698 184315
rect 302187 180980 302253 180981
rect 302187 180916 302188 180980
rect 302252 180916 302253 180980
rect 302187 180915 302253 180916
rect 301635 179076 301701 179077
rect 301635 179012 301636 179076
rect 301700 179012 301701 179076
rect 301635 179011 301701 179012
rect 301635 177580 301701 177581
rect 301635 177516 301636 177580
rect 301700 177516 301701 177580
rect 301635 177515 301701 177516
rect 301638 157861 301698 177515
rect 302190 177309 302250 180915
rect 302187 177308 302253 177309
rect 302187 177244 302188 177308
rect 302252 177244 302253 177308
rect 302187 177243 302253 177244
rect 301819 174588 301885 174589
rect 301819 174524 301820 174588
rect 301884 174524 301885 174588
rect 301819 174523 301885 174524
rect 301635 157860 301701 157861
rect 301635 157796 301636 157860
rect 301700 157796 301701 157860
rect 301635 157795 301701 157796
rect 301822 155549 301882 174523
rect 302374 171150 302434 187990
rect 337147 187938 337189 188174
rect 337425 187938 337467 188174
rect 337147 187854 337467 187938
rect 337147 187618 337189 187854
rect 337425 187618 337467 187854
rect 337147 187586 337467 187618
rect 404744 188174 405064 188206
rect 404744 187938 404786 188174
rect 405022 187938 405064 188174
rect 404744 187854 405064 187938
rect 404744 187618 404786 187854
rect 405022 187618 405064 187854
rect 404744 187586 405064 187618
rect 472341 188174 472661 188206
rect 472341 187938 472383 188174
rect 472619 187938 472661 188174
rect 472341 187854 472661 187938
rect 472341 187618 472383 187854
rect 472619 187618 472661 187854
rect 472341 187586 472661 187618
rect 539938 188174 540258 188206
rect 539938 187938 539980 188174
rect 540216 187938 540258 188174
rect 539938 187854 540258 187938
rect 539938 187618 539980 187854
rect 540216 187618 540258 187854
rect 539938 187586 540258 187618
rect 303349 184454 303669 184486
rect 303349 184218 303391 184454
rect 303627 184218 303669 184454
rect 303349 184134 303669 184218
rect 303349 183898 303391 184134
rect 303627 183898 303669 184134
rect 303349 183866 303669 183898
rect 370946 184454 371266 184486
rect 370946 184218 370988 184454
rect 371224 184218 371266 184454
rect 370946 184134 371266 184218
rect 370946 183898 370988 184134
rect 371224 183898 371266 184134
rect 370946 183866 371266 183898
rect 438543 184454 438863 184486
rect 438543 184218 438585 184454
rect 438821 184218 438863 184454
rect 438543 184134 438863 184218
rect 438543 183898 438585 184134
rect 438821 183898 438863 184134
rect 438543 183866 438863 183898
rect 506140 184454 506460 184486
rect 506140 184218 506182 184454
rect 506418 184218 506460 184454
rect 506140 184134 506460 184218
rect 506140 183898 506182 184134
rect 506418 183898 506460 184134
rect 506140 183866 506460 183898
rect 302555 179892 302621 179893
rect 302555 179828 302556 179892
rect 302620 179890 302621 179892
rect 302620 179830 302802 179890
rect 302620 179828 302621 179830
rect 302555 179827 302621 179828
rect 302374 171090 302618 171150
rect 301819 155548 301885 155549
rect 301819 155484 301820 155548
rect 301884 155484 301885 155548
rect 301819 155483 301885 155484
rect 301454 74490 301698 74550
rect 301083 69188 301149 69189
rect 301083 69124 301084 69188
rect 301148 69124 301149 69188
rect 301083 69123 301149 69124
rect 300163 68916 300229 68917
rect 300163 68852 300164 68916
rect 300228 68852 300229 68916
rect 300163 68851 300229 68852
rect 301086 68781 301146 69123
rect 301638 69053 301698 74490
rect 301635 69052 301701 69053
rect 301635 68988 301636 69052
rect 301700 68988 301701 69052
rect 301635 68987 301701 68988
rect 301083 68780 301149 68781
rect 301083 68716 301084 68780
rect 301148 68716 301149 68780
rect 301083 68715 301149 68716
rect 300347 68644 300413 68645
rect 300347 68580 300348 68644
rect 300412 68580 300413 68644
rect 300347 68579 300413 68580
rect 299979 67964 300045 67965
rect 299979 67900 299980 67964
rect 300044 67900 300045 67964
rect 299979 67899 300045 67900
rect 299795 67556 299861 67557
rect 299795 67492 299796 67556
rect 299860 67492 299861 67556
rect 299795 67491 299861 67492
rect 299611 67012 299677 67013
rect 299611 66948 299612 67012
rect 299676 66948 299677 67012
rect 299611 66947 299677 66948
rect 299614 66605 299674 66947
rect 299611 66604 299677 66605
rect 299611 66540 299612 66604
rect 299676 66540 299677 66604
rect 299611 66539 299677 66540
rect 299614 65620 299674 66539
rect 299982 65620 300042 67899
rect 300350 67829 300410 68579
rect 300531 68508 300597 68509
rect 300531 68444 300532 68508
rect 300596 68444 300597 68508
rect 300531 68443 300597 68444
rect 300347 67828 300413 67829
rect 300347 67764 300348 67828
rect 300412 67764 300413 67828
rect 300347 67763 300413 67764
rect 300350 65620 300410 67763
rect 300534 65925 300594 68443
rect 300531 65924 300597 65925
rect 300531 65860 300532 65924
rect 300596 65860 300597 65924
rect 300531 65859 300597 65860
rect 300534 65650 300594 65859
rect 300534 65590 300748 65650
rect 301086 65620 301146 68715
rect 301451 67556 301517 67557
rect 301451 67492 301452 67556
rect 301516 67492 301517 67556
rect 301451 67491 301517 67492
rect 301454 65620 301514 67491
rect 301638 65650 301698 68987
rect 302187 66876 302253 66877
rect 302187 66812 302188 66876
rect 302252 66812 302253 66876
rect 302187 66811 302253 66812
rect 301638 65590 301852 65650
rect 302190 65620 302250 66811
rect 302558 65620 302618 171090
rect 302742 67557 302802 179830
rect 303294 179830 303600 179890
rect 303107 179212 303173 179213
rect 303107 179148 303108 179212
rect 303172 179148 303173 179212
rect 303107 179147 303173 179148
rect 303110 157317 303170 179147
rect 303294 178870 303354 179830
rect 303294 178810 303600 178870
rect 304306 178840 304366 179520
rect 305042 178840 305102 179520
rect 305778 178500 305838 179520
rect 306514 178840 306574 179520
rect 307250 178840 307310 179520
rect 307986 178840 308046 179520
rect 308722 178840 308782 179520
rect 309458 178840 309518 179520
rect 310194 178840 310254 179520
rect 310930 178840 310990 179520
rect 311666 178876 311726 179520
rect 312402 178876 312462 179520
rect 313138 178876 313198 179520
rect 313874 178876 313934 179520
rect 314610 178876 314670 179520
rect 315346 178876 315406 179520
rect 316082 178876 316142 179520
rect 316818 179430 316878 179520
rect 316818 179370 317154 179430
rect 317094 178870 317154 179370
rect 316848 178810 317154 178870
rect 317554 178840 317614 179520
rect 318290 178840 318350 179520
rect 319026 178840 319086 179520
rect 319762 178840 319822 179520
rect 320498 178840 320558 179520
rect 321234 178500 321294 179520
rect 321970 178840 322030 179520
rect 322706 178840 322766 179520
rect 323442 178840 323502 179520
rect 324178 178840 324238 179520
rect 324914 178840 324974 179520
rect 325650 178840 325710 179520
rect 326386 178840 326446 179520
rect 327122 178840 327182 179520
rect 327858 178840 327918 179520
rect 328594 178840 328654 179520
rect 329330 178840 329390 179520
rect 330066 178840 330126 179520
rect 330802 178840 330862 179520
rect 331538 178840 331598 179520
rect 332274 178840 332334 179520
rect 333010 178840 333070 179520
rect 333746 178840 333806 179520
rect 334482 178840 334542 179520
rect 335123 178940 335189 178941
rect 335123 178876 335124 178940
rect 335188 178876 335189 178940
rect 335123 178875 335189 178876
rect 307365 177879 307685 177936
rect 307365 177643 307407 177879
rect 307643 177643 307685 177879
rect 307365 177586 307685 177643
rect 315207 177879 315527 177936
rect 315207 177643 315249 177879
rect 315485 177643 315527 177879
rect 315207 177586 315527 177643
rect 323049 177879 323369 177936
rect 323049 177643 323091 177879
rect 323327 177643 323369 177879
rect 323049 177586 323369 177643
rect 330891 177879 331211 177936
rect 330891 177643 330933 177879
rect 331169 177643 331211 177879
rect 330891 177586 331211 177643
rect 303444 174454 303764 174486
rect 303444 174218 303486 174454
rect 303722 174218 303764 174454
rect 303444 174134 303764 174218
rect 303444 173898 303486 174134
rect 303722 173898 303764 174134
rect 303444 173866 303764 173898
rect 311286 174454 311606 174486
rect 311286 174218 311328 174454
rect 311564 174218 311606 174454
rect 311286 174134 311606 174218
rect 311286 173898 311328 174134
rect 311564 173898 311606 174134
rect 311286 173866 311606 173898
rect 319128 174454 319448 174486
rect 319128 174218 319170 174454
rect 319406 174218 319448 174454
rect 319128 174134 319448 174218
rect 319128 173898 319170 174134
rect 319406 173898 319448 174134
rect 319128 173866 319448 173898
rect 326970 174454 327290 174486
rect 326970 174218 327012 174454
rect 327248 174218 327290 174454
rect 326970 174134 327290 174218
rect 326970 173898 327012 174134
rect 327248 173898 327290 174134
rect 326970 173866 327290 173898
rect 307365 168174 307685 168206
rect 307365 167938 307407 168174
rect 307643 167938 307685 168174
rect 307365 167854 307685 167938
rect 307365 167618 307407 167854
rect 307643 167618 307685 167854
rect 307365 167586 307685 167618
rect 315207 168174 315527 168206
rect 315207 167938 315249 168174
rect 315485 167938 315527 168174
rect 315207 167854 315527 167938
rect 315207 167618 315249 167854
rect 315485 167618 315527 167854
rect 315207 167586 315527 167618
rect 323049 168174 323369 168206
rect 323049 167938 323091 168174
rect 323327 167938 323369 168174
rect 323049 167854 323369 167938
rect 323049 167618 323091 167854
rect 323327 167618 323369 167854
rect 323049 167586 323369 167618
rect 330891 168174 331211 168206
rect 330891 167938 330933 168174
rect 331169 167938 331211 168174
rect 330891 167854 331211 167938
rect 330891 167618 330933 167854
rect 331169 167618 331211 167854
rect 330891 167586 331211 167618
rect 303444 164454 303764 164486
rect 303444 164218 303486 164454
rect 303722 164218 303764 164454
rect 303444 164134 303764 164218
rect 303444 163898 303486 164134
rect 303722 163898 303764 164134
rect 303444 163866 303764 163898
rect 311286 164454 311606 164486
rect 311286 164218 311328 164454
rect 311564 164218 311606 164454
rect 311286 164134 311606 164218
rect 311286 163898 311328 164134
rect 311564 163898 311606 164134
rect 311286 163866 311606 163898
rect 319128 164454 319448 164486
rect 319128 164218 319170 164454
rect 319406 164218 319448 164454
rect 319128 164134 319448 164218
rect 319128 163898 319170 164134
rect 319406 163898 319448 164134
rect 319128 163866 319448 163898
rect 326970 164454 327290 164486
rect 326970 164218 327012 164454
rect 327248 164218 327290 164454
rect 326970 164134 327290 164218
rect 326970 163898 327012 164134
rect 327248 163898 327290 164134
rect 326970 163866 327290 163898
rect 304947 157996 305013 157997
rect 304947 157932 304948 157996
rect 305012 157932 305013 157996
rect 304947 157931 305013 157932
rect 303107 157316 303173 157317
rect 303107 157252 303108 157316
rect 303172 157252 303173 157316
rect 303107 157251 303173 157252
rect 304395 156772 304461 156773
rect 304395 156708 304396 156772
rect 304460 156708 304461 156772
rect 304395 156707 304461 156708
rect 303475 69596 303541 69597
rect 303475 69532 303476 69596
rect 303540 69532 303541 69596
rect 303475 69531 303541 69532
rect 302739 67556 302805 67557
rect 302739 67492 302740 67556
rect 302804 67492 302805 67556
rect 302739 67491 302805 67492
rect 303478 65620 303538 69531
rect 304398 68917 304458 156707
rect 304950 156637 305010 157931
rect 306051 156908 306117 156909
rect 306051 156844 306052 156908
rect 306116 156844 306117 156908
rect 306051 156843 306117 156844
rect 304947 156636 305013 156637
rect 304947 156572 304948 156636
rect 305012 156572 305013 156636
rect 304947 156571 305013 156572
rect 304211 68916 304277 68917
rect 304211 68852 304212 68916
rect 304276 68852 304277 68916
rect 304211 68851 304277 68852
rect 304395 68916 304461 68917
rect 304395 68852 304396 68916
rect 304460 68852 304461 68916
rect 304395 68851 304461 68852
rect 305683 68916 305749 68917
rect 305683 68852 305684 68916
rect 305748 68852 305749 68916
rect 305683 68851 305749 68852
rect 303843 67556 303909 67557
rect 303843 67492 303844 67556
rect 303908 67492 303909 67556
rect 303843 67491 303909 67492
rect 303846 65620 303906 67491
rect 304214 65620 304274 68851
rect 305315 68372 305381 68373
rect 305315 68308 305316 68372
rect 305380 68308 305381 68372
rect 305315 68307 305381 68308
rect 304579 68236 304645 68237
rect 304579 68172 304580 68236
rect 304644 68172 304645 68236
rect 304579 68171 304645 68172
rect 304582 65620 304642 68171
rect 304947 67556 305013 67557
rect 304947 67492 304948 67556
rect 305012 67492 305013 67556
rect 304947 67491 305013 67492
rect 304950 65620 305010 67491
rect 305318 65620 305378 68307
rect 305686 65620 305746 68851
rect 306054 65620 306114 156843
rect 314699 156636 314765 156637
rect 314699 156572 314700 156636
rect 314764 156572 314765 156636
rect 314699 156571 314765 156572
rect 313227 155548 313293 155549
rect 313227 155484 313228 155548
rect 313292 155484 313293 155548
rect 313227 155483 313293 155484
rect 308627 90404 308693 90405
rect 308627 90340 308628 90404
rect 308692 90340 308693 90404
rect 308627 90339 308693 90340
rect 307155 87548 307221 87549
rect 307155 87484 307156 87548
rect 307220 87484 307221 87548
rect 307155 87483 307221 87484
rect 306419 68916 306485 68917
rect 306419 68852 306420 68916
rect 306484 68852 306485 68916
rect 306419 68851 306485 68852
rect 306422 65620 306482 68851
rect 306787 68236 306853 68237
rect 306787 68172 306788 68236
rect 306852 68172 306853 68236
rect 306787 68171 306853 68172
rect 306790 65620 306850 68171
rect 307158 65620 307218 87483
rect 307523 72452 307589 72453
rect 307523 72388 307524 72452
rect 307588 72388 307589 72452
rect 307523 72387 307589 72388
rect 307526 65620 307586 72387
rect 307891 71092 307957 71093
rect 307891 71028 307892 71092
rect 307956 71028 307957 71092
rect 307891 71027 307957 71028
rect 307894 65620 307954 71027
rect 308259 69596 308325 69597
rect 308259 69532 308260 69596
rect 308324 69532 308325 69596
rect 308259 69531 308325 69532
rect 308262 65620 308322 69531
rect 308630 65620 308690 90339
rect 311019 89044 311085 89045
rect 311019 88980 311020 89044
rect 311084 88980 311085 89044
rect 311019 88979 311085 88980
rect 309363 86188 309429 86189
rect 309363 86124 309364 86188
rect 309428 86124 309429 86188
rect 309363 86123 309429 86124
rect 308995 75172 309061 75173
rect 308995 75108 308996 75172
rect 309060 75108 309061 75172
rect 308995 75107 309061 75108
rect 308998 65620 309058 75107
rect 309366 65620 309426 86123
rect 292992 64171 293312 64240
rect 292992 63935 293034 64171
rect 293270 63935 293312 64171
rect 292992 63866 293312 63935
rect 274035 62796 274101 62797
rect 274035 62732 274036 62796
rect 274100 62732 274101 62796
rect 274035 62731 274101 62732
rect 277632 58174 277952 58206
rect 277632 57938 277674 58174
rect 277910 57938 277952 58174
rect 277632 57854 277952 57938
rect 277632 57618 277674 57854
rect 277910 57618 277952 57854
rect 277632 57586 277952 57618
rect 308352 58174 308672 58206
rect 308352 57938 308394 58174
rect 308630 57938 308672 58174
rect 308352 57854 308672 57938
rect 308352 57618 308394 57854
rect 308630 57618 308672 57854
rect 308352 57586 308672 57618
rect 292992 54454 293312 54486
rect 292992 54218 293034 54454
rect 293270 54218 293312 54454
rect 292992 54134 293312 54218
rect 292992 53898 293034 54134
rect 293270 53898 293312 54134
rect 292992 53866 293312 53898
rect 277632 48174 277952 48206
rect 277632 47938 277674 48174
rect 277910 47938 277952 48174
rect 277632 47854 277952 47938
rect 277632 47618 277674 47854
rect 277910 47618 277952 47854
rect 277632 47586 277952 47618
rect 308352 48174 308672 48206
rect 308352 47938 308394 48174
rect 308630 47938 308672 48174
rect 308352 47854 308672 47938
rect 308352 47618 308394 47854
rect 308630 47618 308672 47854
rect 308352 47586 308672 47618
rect 292992 44454 293312 44486
rect 292992 44218 293034 44454
rect 293270 44218 293312 44454
rect 292992 44134 293312 44218
rect 292992 43898 293034 44134
rect 293270 43898 293312 44134
rect 292992 43866 293312 43898
rect 277632 38174 277952 38206
rect 277632 37938 277674 38174
rect 277910 37938 277952 38174
rect 277632 37854 277952 37938
rect 277632 37618 277674 37854
rect 277910 37618 277952 37854
rect 277632 37586 277952 37618
rect 308352 38174 308672 38206
rect 308352 37938 308394 38174
rect 308630 37938 308672 38174
rect 308352 37854 308672 37938
rect 308352 37618 308394 37854
rect 308630 37618 308672 37854
rect 308352 37586 308672 37618
rect 292992 34454 293312 34486
rect 292992 34218 293034 34454
rect 293270 34218 293312 34454
rect 292992 34134 293312 34218
rect 292992 33898 293034 34134
rect 293270 33898 293312 34134
rect 292992 33866 293312 33898
rect 275326 20501 275386 21760
rect 275694 20637 275754 22100
rect 276092 22070 276306 22130
rect 276246 21725 276306 22070
rect 276614 22070 276828 22130
rect 276614 21861 276674 22070
rect 276611 21860 276677 21861
rect 276611 21796 276612 21860
rect 276676 21796 276677 21860
rect 276611 21795 276677 21796
rect 276243 21724 276309 21725
rect 276243 21660 276244 21724
rect 276308 21660 276309 21724
rect 276243 21659 276309 21660
rect 275691 20636 275757 20637
rect 275691 20572 275692 20636
rect 275756 20572 275757 20636
rect 275691 20571 275757 20572
rect 275323 20500 275389 20501
rect 275323 20436 275324 20500
rect 275388 20436 275389 20500
rect 275323 20435 275389 20436
rect 273851 19276 273917 19277
rect 273851 19212 273852 19276
rect 273916 19212 273917 19276
rect 273851 19211 273917 19212
rect 272379 19140 272445 19141
rect 272379 19076 272380 19140
rect 272444 19076 272445 19140
rect 272379 19075 272445 19076
rect 276430 19005 276490 21760
rect 277166 20365 277226 22100
rect 277564 22070 277778 22130
rect 306268 22070 306482 22130
rect 277718 21997 277778 22070
rect 306422 21997 306482 22070
rect 277715 21996 277781 21997
rect 277715 21932 277716 21996
rect 277780 21932 277781 21996
rect 277715 21931 277781 21932
rect 306419 21996 306485 21997
rect 306419 21932 306420 21996
rect 306484 21932 306485 21996
rect 306419 21931 306485 21932
rect 277163 20364 277229 20365
rect 277163 20300 277164 20364
rect 277228 20300 277229 20364
rect 277163 20299 277229 20300
rect 277902 19413 277962 21760
rect 278270 20229 278330 21760
rect 278267 20228 278333 20229
rect 278267 20164 278268 20228
rect 278332 20164 278333 20228
rect 278267 20163 278333 20164
rect 277899 19412 277965 19413
rect 277899 19348 277900 19412
rect 277964 19348 277965 19412
rect 277899 19347 277965 19348
rect 278638 19277 278698 21760
rect 279006 19549 279066 21760
rect 306606 20637 306666 21760
rect 311022 20637 311082 88979
rect 313230 66877 313290 155483
rect 314702 69733 314762 156571
rect 335126 155277 335186 178875
rect 337702 178840 337762 179520
rect 338438 178500 338498 179520
rect 339174 178840 339234 179520
rect 339910 178840 339970 179520
rect 340646 178840 340706 179520
rect 341382 178840 341442 179520
rect 342118 178840 342178 179520
rect 342854 178840 342914 179520
rect 343590 178840 343650 179520
rect 344326 178840 344386 179520
rect 345062 178840 345122 179520
rect 345798 178840 345858 179520
rect 346534 178840 346594 179520
rect 347270 178840 347330 179520
rect 348006 178840 348066 179520
rect 348742 178876 348802 179520
rect 349478 178876 349538 179520
rect 350214 178876 350274 179520
rect 350950 178876 351010 179520
rect 351686 178500 351746 179860
rect 352422 178500 352482 179520
rect 353158 178840 353218 179520
rect 353894 178840 353954 179860
rect 354630 178500 354690 179520
rect 355366 178840 355426 179520
rect 356102 178840 356162 179860
rect 356838 178500 356898 179520
rect 357574 178840 357634 179860
rect 358310 178840 358370 179860
rect 359046 178840 359106 179520
rect 359782 178840 359842 179860
rect 360518 178500 360578 179520
rect 361254 178840 361314 179520
rect 361990 178840 362050 179520
rect 362726 178840 362786 179860
rect 363462 178840 363522 179860
rect 364198 178840 364258 179860
rect 364934 178840 364994 179520
rect 365670 178840 365730 179520
rect 366406 178840 366466 179520
rect 367142 178840 367202 179520
rect 367878 178840 367938 179520
rect 368614 178840 368674 179520
rect 371834 178876 371894 179520
rect 372570 178840 372630 179520
rect 373306 178840 373366 179520
rect 374042 178840 374102 179520
rect 374778 178840 374838 179520
rect 375514 178840 375574 179520
rect 376250 178840 376310 179520
rect 376986 178840 377046 179520
rect 377722 178840 377782 179520
rect 378458 178840 378518 179520
rect 379194 178840 379254 179520
rect 379930 178876 379990 179520
rect 380666 178876 380726 179520
rect 381402 178876 381462 179520
rect 382138 178876 382198 179520
rect 382874 178876 382934 179520
rect 383610 178876 383670 179520
rect 384346 178840 384406 179520
rect 385082 178840 385142 179520
rect 385818 178840 385878 179520
rect 386554 178840 386614 179520
rect 387290 178840 387350 179520
rect 388026 178840 388086 179520
rect 388762 178840 388822 179520
rect 389498 178840 389558 179520
rect 390234 178840 390294 179520
rect 390970 178840 391030 179520
rect 391706 178840 391766 179520
rect 392442 178840 392502 179520
rect 393178 178840 393238 179520
rect 393914 178840 393974 179520
rect 394650 178840 394710 179520
rect 395386 178840 395446 179520
rect 396122 178840 396182 179520
rect 396858 178840 396918 179520
rect 397594 178840 397654 179520
rect 398330 178840 398390 179520
rect 399066 178840 399126 179520
rect 399802 178840 399862 179520
rect 400538 178840 400598 179520
rect 401274 178840 401334 179520
rect 402010 178840 402070 179520
rect 402746 178840 402806 179520
rect 341497 177879 341817 177936
rect 341497 177643 341539 177879
rect 341775 177643 341817 177879
rect 341497 177586 341817 177643
rect 349339 177879 349659 177936
rect 349339 177643 349381 177879
rect 349617 177643 349659 177879
rect 349339 177586 349659 177643
rect 357181 177879 357501 177936
rect 357181 177643 357223 177879
rect 357459 177643 357501 177879
rect 357181 177586 357501 177643
rect 365023 177879 365343 177936
rect 365023 177643 365065 177879
rect 365301 177643 365343 177879
rect 365023 177586 365343 177643
rect 375629 177879 375949 177936
rect 375629 177643 375671 177879
rect 375907 177643 375949 177879
rect 375629 177586 375949 177643
rect 383471 177879 383791 177936
rect 383471 177643 383513 177879
rect 383749 177643 383791 177879
rect 383471 177586 383791 177643
rect 391313 177879 391633 177936
rect 391313 177643 391355 177879
rect 391591 177643 391633 177879
rect 391313 177586 391633 177643
rect 399155 177879 399475 177936
rect 399155 177643 399197 177879
rect 399433 177643 399475 177879
rect 399155 177586 399475 177643
rect 337576 174454 337896 174486
rect 337576 174218 337618 174454
rect 337854 174218 337896 174454
rect 337576 174134 337896 174218
rect 337576 173898 337618 174134
rect 337854 173898 337896 174134
rect 337576 173866 337896 173898
rect 345418 174454 345738 174486
rect 345418 174218 345460 174454
rect 345696 174218 345738 174454
rect 345418 174134 345738 174218
rect 345418 173898 345460 174134
rect 345696 173898 345738 174134
rect 345418 173866 345738 173898
rect 353260 174454 353580 174486
rect 353260 174218 353302 174454
rect 353538 174218 353580 174454
rect 353260 174134 353580 174218
rect 353260 173898 353302 174134
rect 353538 173898 353580 174134
rect 353260 173866 353580 173898
rect 361102 174454 361422 174486
rect 361102 174218 361144 174454
rect 361380 174218 361422 174454
rect 361102 174134 361422 174218
rect 361102 173898 361144 174134
rect 361380 173898 361422 174134
rect 361102 173866 361422 173898
rect 371708 174454 372028 174486
rect 371708 174218 371750 174454
rect 371986 174218 372028 174454
rect 371708 174134 372028 174218
rect 371708 173898 371750 174134
rect 371986 173898 372028 174134
rect 371708 173866 372028 173898
rect 379550 174454 379870 174486
rect 379550 174218 379592 174454
rect 379828 174218 379870 174454
rect 379550 174134 379870 174218
rect 379550 173898 379592 174134
rect 379828 173898 379870 174134
rect 379550 173866 379870 173898
rect 387392 174454 387712 174486
rect 387392 174218 387434 174454
rect 387670 174218 387712 174454
rect 387392 174134 387712 174218
rect 387392 173898 387434 174134
rect 387670 173898 387712 174134
rect 387392 173866 387712 173898
rect 395234 174454 395554 174486
rect 395234 174218 395276 174454
rect 395512 174218 395554 174454
rect 395234 174134 395554 174218
rect 395234 173898 395276 174134
rect 395512 173898 395554 174134
rect 395234 173866 395554 173898
rect 341497 168174 341817 168206
rect 341497 167938 341539 168174
rect 341775 167938 341817 168174
rect 341497 167854 341817 167938
rect 341497 167618 341539 167854
rect 341775 167618 341817 167854
rect 341497 167586 341817 167618
rect 349339 168174 349659 168206
rect 349339 167938 349381 168174
rect 349617 167938 349659 168174
rect 349339 167854 349659 167938
rect 349339 167618 349381 167854
rect 349617 167618 349659 167854
rect 349339 167586 349659 167618
rect 357181 168174 357501 168206
rect 357181 167938 357223 168174
rect 357459 167938 357501 168174
rect 357181 167854 357501 167938
rect 357181 167618 357223 167854
rect 357459 167618 357501 167854
rect 357181 167586 357501 167618
rect 365023 168174 365343 168206
rect 365023 167938 365065 168174
rect 365301 167938 365343 168174
rect 365023 167854 365343 167938
rect 365023 167618 365065 167854
rect 365301 167618 365343 167854
rect 365023 167586 365343 167618
rect 375629 168174 375949 168206
rect 375629 167938 375671 168174
rect 375907 167938 375949 168174
rect 375629 167854 375949 167938
rect 375629 167618 375671 167854
rect 375907 167618 375949 167854
rect 375629 167586 375949 167618
rect 383471 168174 383791 168206
rect 383471 167938 383513 168174
rect 383749 167938 383791 168174
rect 383471 167854 383791 167938
rect 383471 167618 383513 167854
rect 383749 167618 383791 167854
rect 383471 167586 383791 167618
rect 391313 168174 391633 168206
rect 391313 167938 391355 168174
rect 391591 167938 391633 168174
rect 391313 167854 391633 167938
rect 391313 167618 391355 167854
rect 391591 167618 391633 167854
rect 391313 167586 391633 167618
rect 399155 168174 399475 168206
rect 399155 167938 399197 168174
rect 399433 167938 399475 168174
rect 399155 167854 399475 167938
rect 399155 167618 399197 167854
rect 399433 167618 399475 167854
rect 399155 167586 399475 167618
rect 337576 164454 337896 164486
rect 337576 164218 337618 164454
rect 337854 164218 337896 164454
rect 337576 164134 337896 164218
rect 337576 163898 337618 164134
rect 337854 163898 337896 164134
rect 337576 163866 337896 163898
rect 345418 164454 345738 164486
rect 345418 164218 345460 164454
rect 345696 164218 345738 164454
rect 345418 164134 345738 164218
rect 345418 163898 345460 164134
rect 345696 163898 345738 164134
rect 345418 163866 345738 163898
rect 353260 164454 353580 164486
rect 353260 164218 353302 164454
rect 353538 164218 353580 164454
rect 353260 164134 353580 164218
rect 353260 163898 353302 164134
rect 353538 163898 353580 164134
rect 353260 163866 353580 163898
rect 361102 164454 361422 164486
rect 361102 164218 361144 164454
rect 361380 164218 361422 164454
rect 361102 164134 361422 164218
rect 361102 163898 361144 164134
rect 361380 163898 361422 164134
rect 361102 163866 361422 163898
rect 371708 164454 372028 164486
rect 371708 164218 371750 164454
rect 371986 164218 372028 164454
rect 371708 164134 372028 164218
rect 371708 163898 371750 164134
rect 371986 163898 372028 164134
rect 371708 163866 372028 163898
rect 379550 164454 379870 164486
rect 379550 164218 379592 164454
rect 379828 164218 379870 164454
rect 379550 164134 379870 164218
rect 379550 163898 379592 164134
rect 379828 163898 379870 164134
rect 379550 163866 379870 163898
rect 387392 164454 387712 164486
rect 387392 164218 387434 164454
rect 387670 164218 387712 164454
rect 387392 164134 387712 164218
rect 387392 163898 387434 164134
rect 387670 163898 387712 164134
rect 387392 163866 387712 163898
rect 395234 164454 395554 164486
rect 395234 164218 395276 164454
rect 395512 164218 395554 164454
rect 395234 164134 395554 164218
rect 395234 163898 395276 164134
rect 395512 163898 395554 164134
rect 395234 163866 395554 163898
rect 341497 158174 341817 158206
rect 341497 157938 341539 158174
rect 341775 157938 341817 158174
rect 341497 157854 341817 157938
rect 341497 157618 341539 157854
rect 341775 157618 341817 157854
rect 341497 157586 341817 157618
rect 349339 158174 349659 158206
rect 349339 157938 349381 158174
rect 349617 157938 349659 158174
rect 349339 157854 349659 157938
rect 349339 157618 349381 157854
rect 349617 157618 349659 157854
rect 349339 157586 349659 157618
rect 357181 158174 357501 158206
rect 357181 157938 357223 158174
rect 357459 157938 357501 158174
rect 357181 157854 357501 157938
rect 357181 157618 357223 157854
rect 357459 157618 357501 157854
rect 357181 157586 357501 157618
rect 365023 158174 365343 158206
rect 365023 157938 365065 158174
rect 365301 157938 365343 158174
rect 365023 157854 365343 157938
rect 365023 157618 365065 157854
rect 365301 157618 365343 157854
rect 365023 157586 365343 157618
rect 335123 155276 335189 155277
rect 335123 155212 335124 155276
rect 335188 155212 335189 155276
rect 335123 155211 335189 155212
rect 337576 154454 337896 154486
rect 337576 154218 337618 154454
rect 337854 154218 337896 154454
rect 337576 154134 337896 154218
rect 337576 153898 337618 154134
rect 337854 153898 337896 154134
rect 337576 153866 337896 153898
rect 345418 154454 345738 154486
rect 345418 154218 345460 154454
rect 345696 154218 345738 154454
rect 345418 154134 345738 154218
rect 345418 153898 345460 154134
rect 345696 153898 345738 154134
rect 345418 153866 345738 153898
rect 353260 154454 353580 154486
rect 353260 154218 353302 154454
rect 353538 154218 353580 154454
rect 353260 154134 353580 154218
rect 353260 153898 353302 154134
rect 353538 153898 353580 154134
rect 353260 153866 353580 153898
rect 361102 154454 361422 154486
rect 361102 154218 361144 154454
rect 361380 154218 361422 154454
rect 361102 154134 361422 154218
rect 361102 153898 361144 154134
rect 361380 153898 361422 154134
rect 361102 153866 361422 153898
rect 315803 153780 315869 153781
rect 315803 153716 315804 153780
rect 315868 153716 315869 153780
rect 315803 153715 315869 153716
rect 315806 71229 315866 153715
rect 341497 148174 341817 148206
rect 341497 147938 341539 148174
rect 341775 147938 341817 148174
rect 341497 147854 341817 147938
rect 341497 147618 341539 147854
rect 341775 147618 341817 147854
rect 341497 147586 341817 147618
rect 349339 148174 349659 148206
rect 349339 147938 349381 148174
rect 349617 147938 349659 148174
rect 349339 147854 349659 147938
rect 349339 147618 349381 147854
rect 349617 147618 349659 147854
rect 349339 147586 349659 147618
rect 357181 148174 357501 148206
rect 357181 147938 357223 148174
rect 357459 147938 357501 148174
rect 357181 147854 357501 147938
rect 357181 147618 357223 147854
rect 357459 147618 357501 147854
rect 357181 147586 357501 147618
rect 365023 148174 365343 148206
rect 365023 147938 365065 148174
rect 365301 147938 365343 148174
rect 365023 147854 365343 147938
rect 365023 147618 365065 147854
rect 365301 147618 365343 147854
rect 365023 147586 365343 147618
rect 337576 144454 337896 144486
rect 337576 144218 337618 144454
rect 337854 144218 337896 144454
rect 337576 144134 337896 144218
rect 337576 143898 337618 144134
rect 337854 143898 337896 144134
rect 337576 143866 337896 143898
rect 345418 144454 345738 144486
rect 345418 144218 345460 144454
rect 345696 144218 345738 144454
rect 345418 144134 345738 144218
rect 345418 143898 345460 144134
rect 345696 143898 345738 144134
rect 345418 143866 345738 143898
rect 353260 144454 353580 144486
rect 353260 144218 353302 144454
rect 353538 144218 353580 144454
rect 353260 144134 353580 144218
rect 353260 143898 353302 144134
rect 353538 143898 353580 144134
rect 353260 143866 353580 143898
rect 361102 144454 361422 144486
rect 361102 144218 361144 144454
rect 361380 144218 361422 144454
rect 361102 144134 361422 144218
rect 361102 143898 361144 144134
rect 361380 143898 361422 144134
rect 361102 143866 361422 143898
rect 341497 138174 341817 138206
rect 341497 137938 341539 138174
rect 341775 137938 341817 138174
rect 341497 137854 341817 137938
rect 341497 137618 341539 137854
rect 341775 137618 341817 137854
rect 341497 137586 341817 137618
rect 349339 138174 349659 138206
rect 349339 137938 349381 138174
rect 349617 137938 349659 138174
rect 349339 137854 349659 137938
rect 349339 137618 349381 137854
rect 349617 137618 349659 137854
rect 349339 137586 349659 137618
rect 357181 138174 357501 138206
rect 357181 137938 357223 138174
rect 357459 137938 357501 138174
rect 357181 137854 357501 137938
rect 357181 137618 357223 137854
rect 357459 137618 357501 137854
rect 357181 137586 357501 137618
rect 365023 138174 365343 138206
rect 365023 137938 365065 138174
rect 365301 137938 365343 138174
rect 365023 137854 365343 137938
rect 365023 137618 365065 137854
rect 365301 137618 365343 137854
rect 365023 137586 365343 137618
rect 405966 134842 406026 179520
rect 406702 151830 406762 179520
rect 407438 151830 407498 179520
rect 406702 151770 407130 151830
rect 407438 151770 408050 151830
rect 407070 137730 407130 151770
rect 407070 137670 407314 137730
rect 405966 134782 406548 134842
rect 407254 134300 407314 137670
rect 407990 134640 408050 151770
rect 408174 137730 408234 179520
rect 408910 151830 408970 179520
rect 409646 151830 409706 179520
rect 408910 151770 409522 151830
rect 409646 151770 409890 151830
rect 408174 137670 408786 137730
rect 408726 134640 408786 137670
rect 409462 134640 409522 151770
rect 409830 134842 409890 151770
rect 410382 134842 410442 179520
rect 411118 137050 411178 179520
rect 411118 136990 411362 137050
rect 411302 134842 411362 136990
rect 411854 134842 411914 179520
rect 412590 178870 412650 179520
rect 412406 178810 412650 178870
rect 412406 135690 412466 178810
rect 412406 135630 412834 135690
rect 412774 134842 412834 135630
rect 413326 134842 413386 179520
rect 414062 134842 414122 179520
rect 414798 151830 414858 179520
rect 414798 151770 415410 151830
rect 409830 134782 410228 134842
rect 410382 134782 410964 134842
rect 411302 134782 411700 134842
rect 411854 134782 412436 134842
rect 412774 134782 413172 134842
rect 413326 134782 413908 134842
rect 414062 134782 414644 134842
rect 415350 134812 415410 151770
rect 415534 134842 415594 179520
rect 416270 151830 416330 179520
rect 416270 151770 416698 151830
rect 416638 137730 416698 151770
rect 416638 137670 416882 137730
rect 415534 134782 416116 134842
rect 416822 134812 416882 137670
rect 417006 134842 417066 179520
rect 417742 151830 417802 179520
rect 417742 151770 418170 151830
rect 418110 134842 418170 151770
rect 418478 134842 418538 179860
rect 419214 151830 419274 179520
rect 419214 151770 419458 151830
rect 419398 137050 419458 151770
rect 419398 136990 419642 137050
rect 419582 134842 419642 136990
rect 417006 134782 417588 134842
rect 418110 134782 418324 134842
rect 418478 134782 419060 134842
rect 419582 134782 419796 134842
rect 419950 134788 420010 179860
rect 420686 151830 420746 179860
rect 421422 151830 421482 179860
rect 420686 151770 420930 151830
rect 421422 151770 422034 151830
rect 420870 134788 420930 151770
rect 419950 134728 420532 134788
rect 420870 134728 421268 134788
rect 421974 134640 422034 151770
rect 422158 137730 422218 179520
rect 422158 137670 422770 137730
rect 422710 134690 422770 137670
rect 422894 134788 422954 179520
rect 423630 134788 423690 179520
rect 424366 151830 424426 179520
rect 424366 151770 424978 151830
rect 422894 134728 423476 134788
rect 423630 134728 424212 134788
rect 424918 134640 424978 151770
rect 425102 134788 425162 179520
rect 425838 151830 425898 179860
rect 425838 151770 426450 151830
rect 425102 134728 425684 134788
rect 426390 134690 426450 151770
rect 426574 134788 426634 179520
rect 427310 151830 427370 179520
rect 428046 151830 428106 179520
rect 428782 151830 428842 179520
rect 427310 151770 427738 151830
rect 428046 151770 428658 151830
rect 428782 151770 429210 151830
rect 427678 137730 427738 151770
rect 427678 137670 427922 137730
rect 426574 134728 427156 134788
rect 427862 134758 427922 137670
rect 428598 134640 428658 151770
rect 429150 134788 429210 151770
rect 429518 134788 429578 179860
rect 430254 151830 430314 179860
rect 430254 151770 430498 151830
rect 430438 137050 430498 151770
rect 430438 136990 430682 137050
rect 430622 134788 430682 136990
rect 430990 134788 431050 179520
rect 431726 135270 431786 179520
rect 432462 151830 432522 179520
rect 432462 151770 433074 151830
rect 431726 135210 432154 135270
rect 432094 134788 432154 135210
rect 429150 134728 429364 134788
rect 429518 134728 430100 134788
rect 430622 134728 430836 134788
rect 430990 134728 431572 134788
rect 432094 134728 432308 134788
rect 433014 134690 433074 151770
rect 433198 137050 433258 179520
rect 433198 136990 433442 137050
rect 433382 134788 433442 136990
rect 433934 134788 433994 179520
rect 434670 171150 434730 179860
rect 434670 171090 434914 171150
rect 434854 151830 434914 171090
rect 435406 151830 435466 179520
rect 436142 151830 436202 179520
rect 436878 179210 436938 179520
rect 437062 179490 437490 179550
rect 437062 179210 437122 179490
rect 436878 179150 437122 179210
rect 434854 151770 435282 151830
rect 435406 151770 436018 151830
rect 436142 151770 436754 151830
rect 433382 134728 433780 134788
rect 433934 134728 434516 134788
rect 435222 134640 435282 151770
rect 435958 134640 436018 151770
rect 436694 134640 436754 151770
rect 437430 134640 437490 179490
rect 440098 178876 440158 179520
rect 440834 178840 440894 179520
rect 441570 178840 441630 179520
rect 442306 178840 442366 179520
rect 443042 178876 443102 179520
rect 443778 178876 443838 179520
rect 444514 178876 444574 179520
rect 445250 178876 445310 179520
rect 445986 178876 446046 179520
rect 446722 178876 446782 179520
rect 447458 178876 447518 179520
rect 448194 178876 448254 179520
rect 448930 178876 448990 179520
rect 449666 178876 449726 179520
rect 450402 178876 450462 179520
rect 451138 178876 451198 179520
rect 451874 178876 451934 179520
rect 452610 178876 452670 179520
rect 453346 178876 453406 179520
rect 454082 178840 454142 179520
rect 454818 178840 454878 179520
rect 455554 178840 455614 179520
rect 456290 178500 456350 179520
rect 457026 178840 457086 179520
rect 457762 178840 457822 179520
rect 458498 178840 458558 179520
rect 459234 178840 459294 179520
rect 459970 178840 460030 179520
rect 460706 178840 460766 179520
rect 461442 178840 461502 179520
rect 462178 178840 462238 179520
rect 462914 178840 462974 179520
rect 463650 178840 463710 179520
rect 464386 178840 464446 179520
rect 465122 178840 465182 179520
rect 465858 178840 465918 179520
rect 466594 178840 466654 179520
rect 467330 178840 467390 179520
rect 468066 178840 468126 179520
rect 468802 178840 468862 179520
rect 469538 178840 469598 179520
rect 470274 178840 470334 179520
rect 471010 178840 471070 179520
rect 474230 178876 474290 179860
rect 474966 178500 475026 179520
rect 475702 178840 475762 179520
rect 476438 178840 476498 179520
rect 477174 178840 477234 179860
rect 477910 178840 477970 179860
rect 478646 178876 478706 179520
rect 479382 178876 479442 179860
rect 480118 178876 480178 179520
rect 480854 178876 480914 179860
rect 481590 178876 481650 179520
rect 482326 178876 482386 179520
rect 483062 178876 483122 179520
rect 483798 178876 483858 179520
rect 484534 178876 484594 179520
rect 485270 178876 485330 179520
rect 486006 178876 486066 179520
rect 486742 178876 486802 179520
rect 487478 178876 487538 179520
rect 488214 178840 488274 179520
rect 488950 178840 489010 179520
rect 489686 178840 489746 179520
rect 490422 178840 490482 179520
rect 491158 178840 491218 179520
rect 491894 178840 491954 179520
rect 492630 178840 492690 179520
rect 493366 178840 493426 179520
rect 494102 178840 494162 179520
rect 494838 178840 494898 179520
rect 495574 178840 495634 179520
rect 496310 178840 496370 179520
rect 497046 178840 497106 179520
rect 497782 178840 497842 179520
rect 498518 178840 498578 179520
rect 499254 178840 499314 179520
rect 499990 178840 500050 179520
rect 500726 178840 500786 179520
rect 501462 178840 501522 179520
rect 502198 178840 502258 179520
rect 502934 178840 502994 179520
rect 503670 178840 503730 179520
rect 504406 178840 504466 179520
rect 505142 178840 505202 179520
rect 508362 178876 508422 179520
rect 509098 178840 509158 179520
rect 509834 178840 509894 179520
rect 510570 178876 510630 179520
rect 511306 178876 511366 179520
rect 512042 178840 512102 179520
rect 512778 178876 512838 179520
rect 513514 178876 513574 179520
rect 514250 178876 514310 179520
rect 514986 178876 515046 179520
rect 515722 178840 515782 179520
rect 516458 178876 516518 179520
rect 517194 178876 517254 179520
rect 517930 178876 517990 179520
rect 518666 178876 518726 179520
rect 519402 178876 519462 179520
rect 520138 178876 520198 179520
rect 520874 178876 520934 179520
rect 521610 178876 521670 179520
rect 522346 178840 522406 179520
rect 523082 178500 523142 179520
rect 523818 178840 523878 179520
rect 524554 178840 524614 179520
rect 525290 178840 525350 179520
rect 526026 178840 526086 179520
rect 526762 178840 526822 179520
rect 527498 178840 527558 179520
rect 528234 178840 528294 179520
rect 528970 178840 529030 179520
rect 529706 178840 529766 179520
rect 530442 178840 530502 179520
rect 531178 178840 531238 179520
rect 531914 178840 531974 179520
rect 532650 178840 532710 179520
rect 533386 178840 533446 179520
rect 534122 178840 534182 179520
rect 534858 178840 534918 179520
rect 535594 178840 535654 179520
rect 536330 178840 536390 179520
rect 537066 178840 537126 179520
rect 537802 178840 537862 179520
rect 538538 178840 538598 179520
rect 539274 178840 539334 179520
rect 443893 177879 444213 177936
rect 443893 177643 443935 177879
rect 444171 177643 444213 177879
rect 443893 177586 444213 177643
rect 451735 177879 452055 177936
rect 451735 177643 451777 177879
rect 452013 177643 452055 177879
rect 451735 177586 452055 177643
rect 459577 177879 459897 177936
rect 459577 177643 459619 177879
rect 459855 177643 459897 177879
rect 459577 177586 459897 177643
rect 467419 177879 467739 177936
rect 467419 177643 467461 177879
rect 467697 177643 467739 177879
rect 467419 177586 467739 177643
rect 478025 177879 478345 177936
rect 478025 177643 478067 177879
rect 478303 177643 478345 177879
rect 478025 177586 478345 177643
rect 485867 177879 486187 177936
rect 485867 177643 485909 177879
rect 486145 177643 486187 177879
rect 485867 177586 486187 177643
rect 493709 177879 494029 177936
rect 493709 177643 493751 177879
rect 493987 177643 494029 177879
rect 493709 177586 494029 177643
rect 501551 177879 501871 177936
rect 501551 177643 501593 177879
rect 501829 177643 501871 177879
rect 501551 177586 501871 177643
rect 512157 177879 512477 177936
rect 512157 177643 512199 177879
rect 512435 177643 512477 177879
rect 512157 177586 512477 177643
rect 519999 177879 520319 177936
rect 519999 177643 520041 177879
rect 520277 177643 520319 177879
rect 519999 177586 520319 177643
rect 527841 177879 528161 177936
rect 527841 177643 527883 177879
rect 528119 177643 528161 177879
rect 527841 177586 528161 177643
rect 535683 177879 536003 177936
rect 535683 177643 535725 177879
rect 535961 177643 536003 177879
rect 535683 177586 536003 177643
rect 439972 174454 440292 174486
rect 439972 174218 440014 174454
rect 440250 174218 440292 174454
rect 439972 174134 440292 174218
rect 439972 173898 440014 174134
rect 440250 173898 440292 174134
rect 439972 173866 440292 173898
rect 447814 174454 448134 174486
rect 447814 174218 447856 174454
rect 448092 174218 448134 174454
rect 447814 174134 448134 174218
rect 447814 173898 447856 174134
rect 448092 173898 448134 174134
rect 447814 173866 448134 173898
rect 455656 174454 455976 174486
rect 455656 174218 455698 174454
rect 455934 174218 455976 174454
rect 455656 174134 455976 174218
rect 455656 173898 455698 174134
rect 455934 173898 455976 174134
rect 455656 173866 455976 173898
rect 463498 174454 463818 174486
rect 463498 174218 463540 174454
rect 463776 174218 463818 174454
rect 463498 174134 463818 174218
rect 463498 173898 463540 174134
rect 463776 173898 463818 174134
rect 463498 173866 463818 173898
rect 474104 174454 474424 174486
rect 474104 174218 474146 174454
rect 474382 174218 474424 174454
rect 474104 174134 474424 174218
rect 474104 173898 474146 174134
rect 474382 173898 474424 174134
rect 474104 173866 474424 173898
rect 481946 174454 482266 174486
rect 481946 174218 481988 174454
rect 482224 174218 482266 174454
rect 481946 174134 482266 174218
rect 481946 173898 481988 174134
rect 482224 173898 482266 174134
rect 481946 173866 482266 173898
rect 489788 174454 490108 174486
rect 489788 174218 489830 174454
rect 490066 174218 490108 174454
rect 489788 174134 490108 174218
rect 489788 173898 489830 174134
rect 490066 173898 490108 174134
rect 489788 173866 490108 173898
rect 497630 174454 497950 174486
rect 497630 174218 497672 174454
rect 497908 174218 497950 174454
rect 497630 174134 497950 174218
rect 497630 173898 497672 174134
rect 497908 173898 497950 174134
rect 497630 173866 497950 173898
rect 508236 174454 508556 174486
rect 508236 174218 508278 174454
rect 508514 174218 508556 174454
rect 508236 174134 508556 174218
rect 508236 173898 508278 174134
rect 508514 173898 508556 174134
rect 508236 173866 508556 173898
rect 516078 174454 516398 174486
rect 516078 174218 516120 174454
rect 516356 174218 516398 174454
rect 516078 174134 516398 174218
rect 516078 173898 516120 174134
rect 516356 173898 516398 174134
rect 516078 173866 516398 173898
rect 523920 174454 524240 174486
rect 523920 174218 523962 174454
rect 524198 174218 524240 174454
rect 523920 174134 524240 174218
rect 523920 173898 523962 174134
rect 524198 173898 524240 174134
rect 523920 173866 524240 173898
rect 531762 174454 532082 174486
rect 531762 174218 531804 174454
rect 532040 174218 532082 174454
rect 531762 174134 532082 174218
rect 531762 173898 531804 174134
rect 532040 173898 532082 174134
rect 531762 173866 532082 173898
rect 443893 168174 444213 168206
rect 443893 167938 443935 168174
rect 444171 167938 444213 168174
rect 443893 167854 444213 167938
rect 443893 167618 443935 167854
rect 444171 167618 444213 167854
rect 443893 167586 444213 167618
rect 451735 168174 452055 168206
rect 451735 167938 451777 168174
rect 452013 167938 452055 168174
rect 451735 167854 452055 167938
rect 451735 167618 451777 167854
rect 452013 167618 452055 167854
rect 451735 167586 452055 167618
rect 459577 168174 459897 168206
rect 459577 167938 459619 168174
rect 459855 167938 459897 168174
rect 459577 167854 459897 167938
rect 459577 167618 459619 167854
rect 459855 167618 459897 167854
rect 459577 167586 459897 167618
rect 467419 168174 467739 168206
rect 467419 167938 467461 168174
rect 467697 167938 467739 168174
rect 467419 167854 467739 167938
rect 467419 167618 467461 167854
rect 467697 167618 467739 167854
rect 467419 167586 467739 167618
rect 478025 168174 478345 168206
rect 478025 167938 478067 168174
rect 478303 167938 478345 168174
rect 478025 167854 478345 167938
rect 478025 167618 478067 167854
rect 478303 167618 478345 167854
rect 478025 167586 478345 167618
rect 485867 168174 486187 168206
rect 485867 167938 485909 168174
rect 486145 167938 486187 168174
rect 485867 167854 486187 167938
rect 485867 167618 485909 167854
rect 486145 167618 486187 167854
rect 485867 167586 486187 167618
rect 493709 168174 494029 168206
rect 493709 167938 493751 168174
rect 493987 167938 494029 168174
rect 493709 167854 494029 167938
rect 493709 167618 493751 167854
rect 493987 167618 494029 167854
rect 493709 167586 494029 167618
rect 501551 168174 501871 168206
rect 501551 167938 501593 168174
rect 501829 167938 501871 168174
rect 501551 167854 501871 167938
rect 501551 167618 501593 167854
rect 501829 167618 501871 167854
rect 501551 167586 501871 167618
rect 512157 168174 512477 168206
rect 512157 167938 512199 168174
rect 512435 167938 512477 168174
rect 512157 167854 512477 167938
rect 512157 167618 512199 167854
rect 512435 167618 512477 167854
rect 512157 167586 512477 167618
rect 519999 168174 520319 168206
rect 519999 167938 520041 168174
rect 520277 167938 520319 168174
rect 519999 167854 520319 167938
rect 519999 167618 520041 167854
rect 520277 167618 520319 167854
rect 519999 167586 520319 167618
rect 527841 168174 528161 168206
rect 527841 167938 527883 168174
rect 528119 167938 528161 168174
rect 527841 167854 528161 167938
rect 527841 167618 527883 167854
rect 528119 167618 528161 167854
rect 527841 167586 528161 167618
rect 535683 168174 536003 168206
rect 535683 167938 535725 168174
rect 535961 167938 536003 168174
rect 535683 167854 536003 167938
rect 535683 167618 535725 167854
rect 535961 167618 536003 167854
rect 535683 167586 536003 167618
rect 439972 164454 440292 164486
rect 439972 164218 440014 164454
rect 440250 164218 440292 164454
rect 439972 164134 440292 164218
rect 439972 163898 440014 164134
rect 440250 163898 440292 164134
rect 439972 163866 440292 163898
rect 447814 164454 448134 164486
rect 447814 164218 447856 164454
rect 448092 164218 448134 164454
rect 447814 164134 448134 164218
rect 447814 163898 447856 164134
rect 448092 163898 448134 164134
rect 447814 163866 448134 163898
rect 455656 164454 455976 164486
rect 455656 164218 455698 164454
rect 455934 164218 455976 164454
rect 455656 164134 455976 164218
rect 455656 163898 455698 164134
rect 455934 163898 455976 164134
rect 455656 163866 455976 163898
rect 463498 164454 463818 164486
rect 463498 164218 463540 164454
rect 463776 164218 463818 164454
rect 463498 164134 463818 164218
rect 463498 163898 463540 164134
rect 463776 163898 463818 164134
rect 463498 163866 463818 163898
rect 474104 164454 474424 164486
rect 474104 164218 474146 164454
rect 474382 164218 474424 164454
rect 474104 164134 474424 164218
rect 474104 163898 474146 164134
rect 474382 163898 474424 164134
rect 474104 163866 474424 163898
rect 481946 164454 482266 164486
rect 481946 164218 481988 164454
rect 482224 164218 482266 164454
rect 481946 164134 482266 164218
rect 481946 163898 481988 164134
rect 482224 163898 482266 164134
rect 481946 163866 482266 163898
rect 489788 164454 490108 164486
rect 489788 164218 489830 164454
rect 490066 164218 490108 164454
rect 489788 164134 490108 164218
rect 489788 163898 489830 164134
rect 490066 163898 490108 164134
rect 489788 163866 490108 163898
rect 497630 164454 497950 164486
rect 497630 164218 497672 164454
rect 497908 164218 497950 164454
rect 497630 164134 497950 164218
rect 497630 163898 497672 164134
rect 497908 163898 497950 164134
rect 497630 163866 497950 163898
rect 508236 164454 508556 164486
rect 508236 164218 508278 164454
rect 508514 164218 508556 164454
rect 508236 164134 508556 164218
rect 508236 163898 508278 164134
rect 508514 163898 508556 164134
rect 508236 163866 508556 163898
rect 516078 164454 516398 164486
rect 516078 164218 516120 164454
rect 516356 164218 516398 164454
rect 516078 164134 516398 164218
rect 516078 163898 516120 164134
rect 516356 163898 516398 164134
rect 516078 163866 516398 163898
rect 523920 164454 524240 164486
rect 523920 164218 523962 164454
rect 524198 164218 524240 164454
rect 523920 164134 524240 164218
rect 523920 163898 523962 164134
rect 524198 163898 524240 164134
rect 523920 163866 524240 163898
rect 531762 164454 532082 164486
rect 531762 164218 531804 164454
rect 532040 164218 532082 164454
rect 531762 164134 532082 164218
rect 531762 163898 531804 164134
rect 532040 163898 532082 164134
rect 531762 163866 532082 163898
rect 478025 158174 478345 158206
rect 478025 157938 478067 158174
rect 478303 157938 478345 158174
rect 478025 157854 478345 157938
rect 478025 157618 478067 157854
rect 478303 157618 478345 157854
rect 478025 157586 478345 157618
rect 485867 158174 486187 158206
rect 485867 157938 485909 158174
rect 486145 157938 486187 158174
rect 485867 157854 486187 157938
rect 485867 157618 485909 157854
rect 486145 157618 486187 157854
rect 485867 157586 486187 157618
rect 493709 158174 494029 158206
rect 493709 157938 493751 158174
rect 493987 157938 494029 158174
rect 493709 157854 494029 157938
rect 493709 157618 493751 157854
rect 493987 157618 494029 157854
rect 493709 157586 494029 157618
rect 501551 158174 501871 158206
rect 501551 157938 501593 158174
rect 501829 157938 501871 158174
rect 501551 157854 501871 157938
rect 501551 157618 501593 157854
rect 501829 157618 501871 157854
rect 501551 157586 501871 157618
rect 474104 154454 474424 154486
rect 474104 154218 474146 154454
rect 474382 154218 474424 154454
rect 474104 154134 474424 154218
rect 474104 153898 474146 154134
rect 474382 153898 474424 154134
rect 474104 153866 474424 153898
rect 481946 154454 482266 154486
rect 481946 154218 481988 154454
rect 482224 154218 482266 154454
rect 481946 154134 482266 154218
rect 481946 153898 481988 154134
rect 482224 153898 482266 154134
rect 481946 153866 482266 153898
rect 489788 154454 490108 154486
rect 489788 154218 489830 154454
rect 490066 154218 490108 154454
rect 489788 154134 490108 154218
rect 489788 153898 489830 154134
rect 490066 153898 490108 154134
rect 489788 153866 490108 153898
rect 497630 154454 497950 154486
rect 497630 154218 497672 154454
rect 497908 154218 497950 154454
rect 497630 154134 497950 154218
rect 497630 153898 497672 154134
rect 497908 153898 497950 154134
rect 497630 153866 497950 153898
rect 478025 148174 478345 148206
rect 478025 147938 478067 148174
rect 478303 147938 478345 148174
rect 478025 147854 478345 147938
rect 478025 147618 478067 147854
rect 478303 147618 478345 147854
rect 478025 147586 478345 147618
rect 485867 148174 486187 148206
rect 485867 147938 485909 148174
rect 486145 147938 486187 148174
rect 485867 147854 486187 147938
rect 485867 147618 485909 147854
rect 486145 147618 486187 147854
rect 485867 147586 486187 147618
rect 493709 148174 494029 148206
rect 493709 147938 493751 148174
rect 493987 147938 494029 148174
rect 493709 147854 494029 147938
rect 493709 147618 493751 147854
rect 493987 147618 494029 147854
rect 493709 147586 494029 147618
rect 501551 148174 501871 148206
rect 501551 147938 501593 148174
rect 501829 147938 501871 148174
rect 501551 147854 501871 147938
rect 501551 147618 501593 147854
rect 501829 147618 501871 147854
rect 501551 147586 501871 147618
rect 474104 144454 474424 144486
rect 474104 144218 474146 144454
rect 474382 144218 474424 144454
rect 474104 144134 474424 144218
rect 474104 143898 474146 144134
rect 474382 143898 474424 144134
rect 474104 143866 474424 143898
rect 481946 144454 482266 144486
rect 481946 144218 481988 144454
rect 482224 144218 482266 144454
rect 481946 144134 482266 144218
rect 481946 143898 481988 144134
rect 482224 143898 482266 144134
rect 481946 143866 482266 143898
rect 489788 144454 490108 144486
rect 489788 144218 489830 144454
rect 490066 144218 490108 144454
rect 489788 144134 490108 144218
rect 489788 143898 489830 144134
rect 490066 143898 490108 144134
rect 489788 143866 490108 143898
rect 497630 144454 497950 144486
rect 497630 144218 497672 144454
rect 497908 144218 497950 144454
rect 497630 144134 497950 144218
rect 497630 143898 497672 144134
rect 497908 143898 497950 144134
rect 497630 143866 497950 143898
rect 478025 138174 478345 138206
rect 478025 137938 478067 138174
rect 478303 137938 478345 138174
rect 478025 137854 478345 137938
rect 478025 137618 478067 137854
rect 478303 137618 478345 137854
rect 478025 137586 478345 137618
rect 485867 138174 486187 138206
rect 485867 137938 485909 138174
rect 486145 137938 486187 138174
rect 485867 137854 486187 137938
rect 485867 137618 485909 137854
rect 486145 137618 486187 137854
rect 485867 137586 486187 137618
rect 493709 138174 494029 138206
rect 493709 137938 493751 138174
rect 493987 137938 494029 138174
rect 493709 137854 494029 137938
rect 493709 137618 493751 137854
rect 493987 137618 494029 137854
rect 493709 137586 494029 137618
rect 501551 138174 501871 138206
rect 501551 137938 501593 138174
rect 501829 137938 501871 138174
rect 501551 137854 501871 137938
rect 501551 137618 501593 137854
rect 501829 137618 501871 137854
rect 501551 137586 501871 137618
rect 542494 134842 542554 179520
rect 543230 151830 543290 179520
rect 543966 151830 544026 179520
rect 544702 151830 544762 179520
rect 545438 151830 545498 179520
rect 546174 151830 546234 179520
rect 546910 151830 546970 179520
rect 543230 151770 543658 151830
rect 543966 151770 544578 151830
rect 544702 151770 545130 151830
rect 545438 151770 546050 151830
rect 546174 151770 546418 151830
rect 546910 151770 547522 151830
rect 543598 137730 543658 151770
rect 543598 137670 543842 137730
rect 542494 134782 543076 134842
rect 543782 134795 543842 137670
rect 544518 134640 544578 151770
rect 545070 137730 545130 151770
rect 545070 137670 545314 137730
rect 545254 134758 545314 137670
rect 545990 134640 546050 151770
rect 546358 137730 546418 151770
rect 546358 137670 546786 137730
rect 546726 134640 546786 137670
rect 547462 134758 547522 151770
rect 547646 135270 547706 179860
rect 548382 151830 548442 179520
rect 549118 177170 549178 179520
rect 549118 177110 549730 177170
rect 548382 151770 548994 151830
rect 547646 135210 548258 135270
rect 548198 134640 548258 135210
rect 548934 134758 548994 151770
rect 549670 134640 549730 177110
rect 549854 151830 549914 179860
rect 550590 171150 550650 179520
rect 550590 171090 550834 171150
rect 550774 151830 550834 171090
rect 551326 151830 551386 179520
rect 552062 151830 552122 179860
rect 552798 151830 552858 179520
rect 553534 151830 553594 179520
rect 554270 151830 554330 179520
rect 555006 151830 555066 179520
rect 555742 151830 555802 179860
rect 556478 151830 556538 179520
rect 549854 151770 550466 151830
rect 550774 151770 551202 151830
rect 551326 151770 551938 151830
rect 552062 151770 552674 151830
rect 552798 151770 553410 151830
rect 553534 151770 554146 151830
rect 554270 151770 554698 151830
rect 555006 151770 555618 151830
rect 555742 151770 556170 151830
rect 556478 151770 557090 151830
rect 550406 134640 550466 151770
rect 551142 134690 551202 151770
rect 551878 134640 551938 151770
rect 552614 134640 552674 151770
rect 553350 134640 553410 151770
rect 554086 134640 554146 151770
rect 554638 138030 554698 151770
rect 554638 137970 554882 138030
rect 554822 134758 554882 137970
rect 555558 134758 555618 151770
rect 556110 138030 556170 151770
rect 556110 137970 556354 138030
rect 556294 134758 556354 137970
rect 557030 134690 557090 151770
rect 557214 138030 557274 179520
rect 557950 151830 558010 179520
rect 558686 177170 558746 179520
rect 558686 177110 559298 177170
rect 557950 151770 558562 151830
rect 557214 137970 557826 138030
rect 557766 134690 557826 137970
rect 558502 134758 558562 151770
rect 559238 134758 559298 177110
rect 559422 151830 559482 179520
rect 560158 177170 560218 179520
rect 560158 177110 560770 177170
rect 559422 151770 560034 151830
rect 559974 134758 560034 151770
rect 560710 134758 560770 177110
rect 560894 151830 560954 179520
rect 561630 151830 561690 179520
rect 562366 151830 562426 179520
rect 563102 151830 563162 179520
rect 563838 151830 563898 179520
rect 564574 151830 564634 179520
rect 560894 151770 561506 151830
rect 561630 151770 562242 151830
rect 562366 151770 562978 151830
rect 563102 151770 563714 151830
rect 563838 151770 564450 151830
rect 564574 151770 565186 151830
rect 561446 134758 561506 151770
rect 562182 134690 562242 151770
rect 562918 134758 562978 151770
rect 563654 134758 563714 151770
rect 564390 134758 564450 151770
rect 565126 134758 565186 151770
rect 565310 138030 565370 179520
rect 566046 151830 566106 179520
rect 566782 151830 566842 179520
rect 567518 151830 567578 179520
rect 566046 151770 566658 151830
rect 566782 151770 567026 151830
rect 567518 151770 568130 151830
rect 565310 137970 565922 138030
rect 565862 134640 565922 137970
rect 566598 134640 566658 151770
rect 566966 135270 567026 151770
rect 566966 135210 567394 135270
rect 567334 134758 567394 135210
rect 568070 134690 568130 151770
rect 568254 137730 568314 179520
rect 568990 151830 569050 179520
rect 568990 151770 569602 151830
rect 568254 137670 568866 137730
rect 568806 134640 568866 137670
rect 569542 134640 569602 151770
rect 569726 137730 569786 179520
rect 570462 151830 570522 179520
rect 570462 151770 571074 151830
rect 569726 137670 570338 137730
rect 570278 134640 570338 137670
rect 571014 134640 571074 151770
rect 571198 137730 571258 179520
rect 571934 151830 571994 179520
rect 572670 151830 572730 179520
rect 573406 151830 573466 179520
rect 571934 151770 572546 151830
rect 572670 151770 573282 151830
rect 573406 151770 574018 151830
rect 571198 137670 571810 137730
rect 571750 134640 571810 137670
rect 572486 134758 572546 151770
rect 573222 134640 573282 151770
rect 573958 134758 574018 151770
rect 373056 128174 373376 128206
rect 373056 127938 373098 128174
rect 373334 127938 373376 128174
rect 373056 127854 373376 127938
rect 373056 127618 373098 127854
rect 373334 127618 373376 127854
rect 373056 127586 373376 127618
rect 403776 128174 404096 128206
rect 403776 127938 403818 128174
rect 404054 127938 404096 128174
rect 403776 127854 404096 127938
rect 403776 127618 403818 127854
rect 404054 127618 404096 127854
rect 403776 127586 404096 127618
rect 434496 128174 434816 128206
rect 434496 127938 434538 128174
rect 434774 127938 434816 128174
rect 434496 127854 434816 127938
rect 434496 127618 434538 127854
rect 434774 127618 434816 127854
rect 434496 127586 434816 127618
rect 448144 128174 448464 128206
rect 448144 127938 448186 128174
rect 448422 127938 448464 128174
rect 448144 127854 448464 127938
rect 448144 127618 448186 127854
rect 448422 127618 448464 127854
rect 448144 127586 448464 127618
rect 478864 128174 479184 128206
rect 478864 127938 478906 128174
rect 479142 127938 479184 128174
rect 478864 127854 479184 127938
rect 478864 127618 478906 127854
rect 479142 127618 479184 127854
rect 478864 127586 479184 127618
rect 509584 128174 509904 128206
rect 509584 127938 509626 128174
rect 509862 127938 509904 128174
rect 509584 127854 509904 127938
rect 509584 127618 509626 127854
rect 509862 127618 509904 127854
rect 509584 127586 509904 127618
rect 540304 128174 540624 128206
rect 540304 127938 540346 128174
rect 540582 127938 540624 128174
rect 540304 127854 540624 127938
rect 540304 127618 540346 127854
rect 540582 127618 540624 127854
rect 540304 127586 540624 127618
rect 571024 128174 571344 128206
rect 571024 127938 571066 128174
rect 571302 127938 571344 128174
rect 571024 127854 571344 127938
rect 571024 127618 571066 127854
rect 571302 127618 571344 127854
rect 571024 127586 571344 127618
rect 388416 124454 388736 124486
rect 388416 124218 388458 124454
rect 388694 124218 388736 124454
rect 388416 124134 388736 124218
rect 388416 123898 388458 124134
rect 388694 123898 388736 124134
rect 388416 123866 388736 123898
rect 419136 124454 419456 124486
rect 419136 124218 419178 124454
rect 419414 124218 419456 124454
rect 419136 124134 419456 124218
rect 419136 123898 419178 124134
rect 419414 123898 419456 124134
rect 419136 123866 419456 123898
rect 463504 124454 463824 124486
rect 463504 124218 463546 124454
rect 463782 124218 463824 124454
rect 463504 124134 463824 124218
rect 463504 123898 463546 124134
rect 463782 123898 463824 124134
rect 463504 123866 463824 123898
rect 494224 124454 494544 124486
rect 494224 124218 494266 124454
rect 494502 124218 494544 124454
rect 494224 124134 494544 124218
rect 494224 123898 494266 124134
rect 494502 123898 494544 124134
rect 494224 123866 494544 123898
rect 524944 124454 525264 124486
rect 524944 124218 524986 124454
rect 525222 124218 525264 124454
rect 524944 124134 525264 124218
rect 524944 123898 524986 124134
rect 525222 123898 525264 124134
rect 524944 123866 525264 123898
rect 555664 124454 555984 124486
rect 555664 124218 555706 124454
rect 555942 124218 555984 124454
rect 555664 124134 555984 124218
rect 555664 123898 555706 124134
rect 555942 123898 555984 124134
rect 555664 123866 555984 123898
rect 373056 118174 373376 118206
rect 373056 117938 373098 118174
rect 373334 117938 373376 118174
rect 373056 117854 373376 117938
rect 373056 117618 373098 117854
rect 373334 117618 373376 117854
rect 373056 117586 373376 117618
rect 403776 118174 404096 118206
rect 403776 117938 403818 118174
rect 404054 117938 404096 118174
rect 403776 117854 404096 117938
rect 403776 117618 403818 117854
rect 404054 117618 404096 117854
rect 403776 117586 404096 117618
rect 434496 118174 434816 118206
rect 434496 117938 434538 118174
rect 434774 117938 434816 118174
rect 434496 117854 434816 117938
rect 434496 117618 434538 117854
rect 434774 117618 434816 117854
rect 434496 117586 434816 117618
rect 448144 118174 448464 118206
rect 448144 117938 448186 118174
rect 448422 117938 448464 118174
rect 448144 117854 448464 117938
rect 448144 117618 448186 117854
rect 448422 117618 448464 117854
rect 448144 117586 448464 117618
rect 478864 118174 479184 118206
rect 478864 117938 478906 118174
rect 479142 117938 479184 118174
rect 478864 117854 479184 117938
rect 478864 117618 478906 117854
rect 479142 117618 479184 117854
rect 478864 117586 479184 117618
rect 509584 118174 509904 118206
rect 509584 117938 509626 118174
rect 509862 117938 509904 118174
rect 509584 117854 509904 117938
rect 509584 117618 509626 117854
rect 509862 117618 509904 117854
rect 509584 117586 509904 117618
rect 540304 118174 540624 118206
rect 540304 117938 540346 118174
rect 540582 117938 540624 118174
rect 540304 117854 540624 117938
rect 540304 117618 540346 117854
rect 540582 117618 540624 117854
rect 540304 117586 540624 117618
rect 571024 118174 571344 118206
rect 571024 117938 571066 118174
rect 571302 117938 571344 118174
rect 571024 117854 571344 117938
rect 571024 117618 571066 117854
rect 571302 117618 571344 117854
rect 571024 117586 571344 117618
rect 388416 114454 388736 114486
rect 388416 114218 388458 114454
rect 388694 114218 388736 114454
rect 388416 114134 388736 114218
rect 388416 113898 388458 114134
rect 388694 113898 388736 114134
rect 388416 113866 388736 113898
rect 419136 114454 419456 114486
rect 419136 114218 419178 114454
rect 419414 114218 419456 114454
rect 419136 114134 419456 114218
rect 419136 113898 419178 114134
rect 419414 113898 419456 114134
rect 419136 113866 419456 113898
rect 463504 114454 463824 114486
rect 463504 114218 463546 114454
rect 463782 114218 463824 114454
rect 463504 114134 463824 114218
rect 463504 113898 463546 114134
rect 463782 113898 463824 114134
rect 463504 113866 463824 113898
rect 494224 114454 494544 114486
rect 494224 114218 494266 114454
rect 494502 114218 494544 114454
rect 494224 114134 494544 114218
rect 494224 113898 494266 114134
rect 494502 113898 494544 114134
rect 494224 113866 494544 113898
rect 524944 114454 525264 114486
rect 524944 114218 524986 114454
rect 525222 114218 525264 114454
rect 524944 114134 525264 114218
rect 524944 113898 524986 114134
rect 525222 113898 525264 114134
rect 524944 113866 525264 113898
rect 555664 114454 555984 114486
rect 555664 114218 555706 114454
rect 555942 114218 555984 114454
rect 555664 114134 555984 114218
rect 555664 113898 555706 114134
rect 555942 113898 555984 114134
rect 555664 113866 555984 113898
rect 373056 108174 373376 108206
rect 373056 107938 373098 108174
rect 373334 107938 373376 108174
rect 373056 107854 373376 107938
rect 373056 107618 373098 107854
rect 373334 107618 373376 107854
rect 373056 107586 373376 107618
rect 403776 108174 404096 108206
rect 403776 107938 403818 108174
rect 404054 107938 404096 108174
rect 403776 107854 404096 107938
rect 403776 107618 403818 107854
rect 404054 107618 404096 107854
rect 403776 107586 404096 107618
rect 434496 108174 434816 108206
rect 434496 107938 434538 108174
rect 434774 107938 434816 108174
rect 434496 107854 434816 107938
rect 434496 107618 434538 107854
rect 434774 107618 434816 107854
rect 434496 107586 434816 107618
rect 448144 108174 448464 108206
rect 448144 107938 448186 108174
rect 448422 107938 448464 108174
rect 448144 107854 448464 107938
rect 448144 107618 448186 107854
rect 448422 107618 448464 107854
rect 448144 107586 448464 107618
rect 478864 108174 479184 108206
rect 478864 107938 478906 108174
rect 479142 107938 479184 108174
rect 478864 107854 479184 107938
rect 478864 107618 478906 107854
rect 479142 107618 479184 107854
rect 478864 107586 479184 107618
rect 509584 108174 509904 108206
rect 509584 107938 509626 108174
rect 509862 107938 509904 108174
rect 509584 107854 509904 107938
rect 509584 107618 509626 107854
rect 509862 107618 509904 107854
rect 509584 107586 509904 107618
rect 540304 108174 540624 108206
rect 540304 107938 540346 108174
rect 540582 107938 540624 108174
rect 540304 107854 540624 107938
rect 540304 107618 540346 107854
rect 540582 107618 540624 107854
rect 540304 107586 540624 107618
rect 571024 108174 571344 108206
rect 571024 107938 571066 108174
rect 571302 107938 571344 108174
rect 571024 107854 571344 107938
rect 571024 107618 571066 107854
rect 571302 107618 571344 107854
rect 571024 107586 571344 107618
rect 388416 104454 388736 104486
rect 388416 104218 388458 104454
rect 388694 104218 388736 104454
rect 388416 104134 388736 104218
rect 388416 103898 388458 104134
rect 388694 103898 388736 104134
rect 388416 103866 388736 103898
rect 419136 104454 419456 104486
rect 419136 104218 419178 104454
rect 419414 104218 419456 104454
rect 419136 104134 419456 104218
rect 419136 103898 419178 104134
rect 419414 103898 419456 104134
rect 419136 103866 419456 103898
rect 463504 104454 463824 104486
rect 463504 104218 463546 104454
rect 463782 104218 463824 104454
rect 463504 104134 463824 104218
rect 463504 103898 463546 104134
rect 463782 103898 463824 104134
rect 463504 103866 463824 103898
rect 494224 104454 494544 104486
rect 494224 104218 494266 104454
rect 494502 104218 494544 104454
rect 494224 104134 494544 104218
rect 494224 103898 494266 104134
rect 494502 103898 494544 104134
rect 494224 103866 494544 103898
rect 524944 104454 525264 104486
rect 524944 104218 524986 104454
rect 525222 104218 525264 104454
rect 524944 104134 525264 104218
rect 524944 103898 524986 104134
rect 525222 103898 525264 104134
rect 524944 103866 525264 103898
rect 555664 104454 555984 104486
rect 555664 104218 555706 104454
rect 555942 104218 555984 104454
rect 555664 104134 555984 104218
rect 555664 103898 555706 104134
rect 555942 103898 555984 104134
rect 555664 103866 555984 103898
rect 373056 98174 373376 98206
rect 373056 97938 373098 98174
rect 373334 97938 373376 98174
rect 373056 97854 373376 97938
rect 373056 97618 373098 97854
rect 373334 97618 373376 97854
rect 373056 97586 373376 97618
rect 403776 98174 404096 98206
rect 403776 97938 403818 98174
rect 404054 97938 404096 98174
rect 403776 97854 404096 97938
rect 403776 97618 403818 97854
rect 404054 97618 404096 97854
rect 403776 97586 404096 97618
rect 434496 98174 434816 98206
rect 434496 97938 434538 98174
rect 434774 97938 434816 98174
rect 434496 97854 434816 97938
rect 434496 97618 434538 97854
rect 434774 97618 434816 97854
rect 434496 97586 434816 97618
rect 448144 98174 448464 98206
rect 448144 97938 448186 98174
rect 448422 97938 448464 98174
rect 448144 97854 448464 97938
rect 448144 97618 448186 97854
rect 448422 97618 448464 97854
rect 448144 97586 448464 97618
rect 478864 98174 479184 98206
rect 478864 97938 478906 98174
rect 479142 97938 479184 98174
rect 478864 97854 479184 97938
rect 478864 97618 478906 97854
rect 479142 97618 479184 97854
rect 478864 97586 479184 97618
rect 509584 98174 509904 98206
rect 509584 97938 509626 98174
rect 509862 97938 509904 98174
rect 509584 97854 509904 97938
rect 509584 97618 509626 97854
rect 509862 97618 509904 97854
rect 509584 97586 509904 97618
rect 540304 98174 540624 98206
rect 540304 97938 540346 98174
rect 540582 97938 540624 98174
rect 540304 97854 540624 97938
rect 540304 97618 540346 97854
rect 540582 97618 540624 97854
rect 540304 97586 540624 97618
rect 571024 98174 571344 98206
rect 571024 97938 571066 98174
rect 571302 97938 571344 98174
rect 571024 97854 571344 97938
rect 571024 97618 571066 97854
rect 571302 97618 571344 97854
rect 571024 97586 571344 97618
rect 388416 94454 388736 94486
rect 388416 94218 388458 94454
rect 388694 94218 388736 94454
rect 388416 94134 388736 94218
rect 388416 93898 388458 94134
rect 388694 93898 388736 94134
rect 388416 93866 388736 93898
rect 419136 94454 419456 94486
rect 419136 94218 419178 94454
rect 419414 94218 419456 94454
rect 419136 94134 419456 94218
rect 419136 93898 419178 94134
rect 419414 93898 419456 94134
rect 419136 93866 419456 93898
rect 463504 94454 463824 94486
rect 463504 94218 463546 94454
rect 463782 94218 463824 94454
rect 463504 94134 463824 94218
rect 463504 93898 463546 94134
rect 463782 93898 463824 94134
rect 463504 93866 463824 93898
rect 494224 94454 494544 94486
rect 494224 94218 494266 94454
rect 494502 94218 494544 94454
rect 494224 94134 494544 94218
rect 494224 93898 494266 94134
rect 494502 93898 494544 94134
rect 494224 93866 494544 93898
rect 524944 94454 525264 94486
rect 524944 94218 524986 94454
rect 525222 94218 525264 94454
rect 524944 94134 525264 94218
rect 524944 93898 524986 94134
rect 525222 93898 525264 94134
rect 524944 93866 525264 93898
rect 555664 94454 555984 94486
rect 555664 94218 555706 94454
rect 555942 94218 555984 94454
rect 555664 94134 555984 94218
rect 555664 93898 555706 94134
rect 555942 93898 555984 94134
rect 555664 93866 555984 93898
rect 315803 71228 315869 71229
rect 315803 71164 315804 71228
rect 315868 71164 315869 71228
rect 315803 71163 315869 71164
rect 574694 71093 574754 564299
rect 574875 511324 574941 511325
rect 574875 511260 574876 511324
rect 574940 511260 574941 511324
rect 574875 511259 574941 511260
rect 574691 71092 574757 71093
rect 574691 71028 574692 71092
rect 574756 71028 574757 71092
rect 574691 71027 574757 71028
rect 314699 69732 314765 69733
rect 314699 69668 314700 69732
rect 314764 69668 314765 69732
rect 314699 69667 314765 69668
rect 574878 69597 574938 511259
rect 575982 87549 576042 670651
rect 585310 668174 585930 677618
rect 585310 667938 585342 668174
rect 585578 667938 585662 668174
rect 585898 667938 585930 668174
rect 585310 667854 585930 667938
rect 585310 667618 585342 667854
rect 585578 667618 585662 667854
rect 585898 667618 585930 667854
rect 585310 658174 585930 667618
rect 585310 657938 585342 658174
rect 585578 657938 585662 658174
rect 585898 657938 585930 658174
rect 585310 657854 585930 657938
rect 585310 657618 585342 657854
rect 585578 657618 585662 657854
rect 585898 657618 585930 657854
rect 585310 648174 585930 657618
rect 585310 647938 585342 648174
rect 585578 647938 585662 648174
rect 585898 647938 585930 648174
rect 585310 647854 585930 647938
rect 585310 647618 585342 647854
rect 585578 647618 585662 647854
rect 585898 647618 585930 647854
rect 585310 638174 585930 647618
rect 585310 637938 585342 638174
rect 585578 637938 585662 638174
rect 585898 637938 585930 638174
rect 585310 637854 585930 637938
rect 585310 637618 585342 637854
rect 585578 637618 585662 637854
rect 585898 637618 585930 637854
rect 585310 628174 585930 637618
rect 585310 627938 585342 628174
rect 585578 627938 585662 628174
rect 585898 627938 585930 628174
rect 585310 627854 585930 627938
rect 585310 627618 585342 627854
rect 585578 627618 585662 627854
rect 585898 627618 585930 627854
rect 585310 618174 585930 627618
rect 585310 617938 585342 618174
rect 585578 617938 585662 618174
rect 585898 617938 585930 618174
rect 585310 617854 585930 617938
rect 585310 617618 585342 617854
rect 585578 617618 585662 617854
rect 585898 617618 585930 617854
rect 576163 617540 576229 617541
rect 576163 617476 576164 617540
rect 576228 617476 576229 617540
rect 576163 617475 576229 617476
rect 575979 87548 576045 87549
rect 575979 87484 575980 87548
rect 576044 87484 576045 87548
rect 575979 87483 576045 87484
rect 576166 72453 576226 617475
rect 585310 608174 585930 617618
rect 585310 607938 585342 608174
rect 585578 607938 585662 608174
rect 585898 607938 585930 608174
rect 585310 607854 585930 607938
rect 585310 607618 585342 607854
rect 585578 607618 585662 607854
rect 585898 607618 585930 607854
rect 585310 598174 585930 607618
rect 585310 597938 585342 598174
rect 585578 597938 585662 598174
rect 585898 597938 585930 598174
rect 585310 597854 585930 597938
rect 585310 597618 585342 597854
rect 585578 597618 585662 597854
rect 585898 597618 585930 597854
rect 585310 588174 585930 597618
rect 585310 587938 585342 588174
rect 585578 587938 585662 588174
rect 585898 587938 585930 588174
rect 585310 587854 585930 587938
rect 585310 587618 585342 587854
rect 585578 587618 585662 587854
rect 585898 587618 585930 587854
rect 585310 578174 585930 587618
rect 585310 577938 585342 578174
rect 585578 577938 585662 578174
rect 585898 577938 585930 578174
rect 585310 577854 585930 577938
rect 585310 577618 585342 577854
rect 585578 577618 585662 577854
rect 585898 577618 585930 577854
rect 585310 568174 585930 577618
rect 585310 567938 585342 568174
rect 585578 567938 585662 568174
rect 585898 567938 585930 568174
rect 585310 567854 585930 567938
rect 585310 567618 585342 567854
rect 585578 567618 585662 567854
rect 585898 567618 585930 567854
rect 585310 558174 585930 567618
rect 585310 557938 585342 558174
rect 585578 557938 585662 558174
rect 585898 557938 585930 558174
rect 585310 557854 585930 557938
rect 585310 557618 585342 557854
rect 585578 557618 585662 557854
rect 585898 557618 585930 557854
rect 585310 548174 585930 557618
rect 585310 547938 585342 548174
rect 585578 547938 585662 548174
rect 585898 547938 585930 548174
rect 585310 547854 585930 547938
rect 585310 547618 585342 547854
rect 585578 547618 585662 547854
rect 585898 547618 585930 547854
rect 585310 538174 585930 547618
rect 585310 537938 585342 538174
rect 585578 537938 585662 538174
rect 585898 537938 585930 538174
rect 585310 537854 585930 537938
rect 585310 537618 585342 537854
rect 585578 537618 585662 537854
rect 585898 537618 585930 537854
rect 585310 528174 585930 537618
rect 585310 527938 585342 528174
rect 585578 527938 585662 528174
rect 585898 527938 585930 528174
rect 585310 527854 585930 527938
rect 585310 527618 585342 527854
rect 585578 527618 585662 527854
rect 585898 527618 585930 527854
rect 585310 518174 585930 527618
rect 585310 517938 585342 518174
rect 585578 517938 585662 518174
rect 585898 517938 585930 518174
rect 585310 517854 585930 517938
rect 585310 517618 585342 517854
rect 585578 517618 585662 517854
rect 585898 517618 585930 517854
rect 585310 508174 585930 517618
rect 585310 507938 585342 508174
rect 585578 507938 585662 508174
rect 585898 507938 585930 508174
rect 585310 507854 585930 507938
rect 585310 507618 585342 507854
rect 585578 507618 585662 507854
rect 585898 507618 585930 507854
rect 585310 498174 585930 507618
rect 585310 497938 585342 498174
rect 585578 497938 585662 498174
rect 585898 497938 585930 498174
rect 585310 497854 585930 497938
rect 585310 497618 585342 497854
rect 585578 497618 585662 497854
rect 585898 497618 585930 497854
rect 585310 488174 585930 497618
rect 585310 487938 585342 488174
rect 585578 487938 585662 488174
rect 585898 487938 585930 488174
rect 585310 487854 585930 487938
rect 585310 487618 585342 487854
rect 585578 487618 585662 487854
rect 585898 487618 585930 487854
rect 585310 478174 585930 487618
rect 585310 477938 585342 478174
rect 585578 477938 585662 478174
rect 585898 477938 585930 478174
rect 585310 477854 585930 477938
rect 585310 477618 585342 477854
rect 585578 477618 585662 477854
rect 585898 477618 585930 477854
rect 585310 468174 585930 477618
rect 585310 467938 585342 468174
rect 585578 467938 585662 468174
rect 585898 467938 585930 468174
rect 585310 467854 585930 467938
rect 585310 467618 585342 467854
rect 585578 467618 585662 467854
rect 585898 467618 585930 467854
rect 585310 458174 585930 467618
rect 578739 458148 578805 458149
rect 578739 458084 578740 458148
rect 578804 458084 578805 458148
rect 578739 458083 578805 458084
rect 577451 404972 577517 404973
rect 577451 404908 577452 404972
rect 577516 404908 577517 404972
rect 577451 404907 577517 404908
rect 577454 75173 577514 404907
rect 577635 351932 577701 351933
rect 577635 351868 577636 351932
rect 577700 351868 577701 351932
rect 577635 351867 577701 351868
rect 577638 86189 577698 351867
rect 578742 90405 578802 458083
rect 585310 457938 585342 458174
rect 585578 457938 585662 458174
rect 585898 457938 585930 458174
rect 585310 457854 585930 457938
rect 585310 457618 585342 457854
rect 585578 457618 585662 457854
rect 585898 457618 585930 457854
rect 585310 448174 585930 457618
rect 585310 447938 585342 448174
rect 585578 447938 585662 448174
rect 585898 447938 585930 448174
rect 585310 447854 585930 447938
rect 585310 447618 585342 447854
rect 585578 447618 585662 447854
rect 585898 447618 585930 447854
rect 585310 438174 585930 447618
rect 585310 437938 585342 438174
rect 585578 437938 585662 438174
rect 585898 437938 585930 438174
rect 585310 437854 585930 437938
rect 585310 437618 585342 437854
rect 585578 437618 585662 437854
rect 585898 437618 585930 437854
rect 585310 428174 585930 437618
rect 585310 427938 585342 428174
rect 585578 427938 585662 428174
rect 585898 427938 585930 428174
rect 585310 427854 585930 427938
rect 585310 427618 585342 427854
rect 585578 427618 585662 427854
rect 585898 427618 585930 427854
rect 585310 418174 585930 427618
rect 585310 417938 585342 418174
rect 585578 417938 585662 418174
rect 585898 417938 585930 418174
rect 585310 417854 585930 417938
rect 585310 417618 585342 417854
rect 585578 417618 585662 417854
rect 585898 417618 585930 417854
rect 585310 408174 585930 417618
rect 585310 407938 585342 408174
rect 585578 407938 585662 408174
rect 585898 407938 585930 408174
rect 585310 407854 585930 407938
rect 585310 407618 585342 407854
rect 585578 407618 585662 407854
rect 585898 407618 585930 407854
rect 585310 398174 585930 407618
rect 585310 397938 585342 398174
rect 585578 397938 585662 398174
rect 585898 397938 585930 398174
rect 585310 397854 585930 397938
rect 585310 397618 585342 397854
rect 585578 397618 585662 397854
rect 585898 397618 585930 397854
rect 585310 388174 585930 397618
rect 585310 387938 585342 388174
rect 585578 387938 585662 388174
rect 585898 387938 585930 388174
rect 585310 387854 585930 387938
rect 585310 387618 585342 387854
rect 585578 387618 585662 387854
rect 585898 387618 585930 387854
rect 585310 378174 585930 387618
rect 585310 377938 585342 378174
rect 585578 377938 585662 378174
rect 585898 377938 585930 378174
rect 585310 377854 585930 377938
rect 585310 377618 585342 377854
rect 585578 377618 585662 377854
rect 585898 377618 585930 377854
rect 585310 368174 585930 377618
rect 585310 367938 585342 368174
rect 585578 367938 585662 368174
rect 585898 367938 585930 368174
rect 585310 367854 585930 367938
rect 585310 367618 585342 367854
rect 585578 367618 585662 367854
rect 585898 367618 585930 367854
rect 585310 358174 585930 367618
rect 585310 357938 585342 358174
rect 585578 357938 585662 358174
rect 585898 357938 585930 358174
rect 585310 357854 585930 357938
rect 585310 357618 585342 357854
rect 585578 357618 585662 357854
rect 585898 357618 585930 357854
rect 585310 348174 585930 357618
rect 585310 347938 585342 348174
rect 585578 347938 585662 348174
rect 585898 347938 585930 348174
rect 585310 347854 585930 347938
rect 585310 347618 585342 347854
rect 585578 347618 585662 347854
rect 585898 347618 585930 347854
rect 585310 338174 585930 347618
rect 585310 337938 585342 338174
rect 585578 337938 585662 338174
rect 585898 337938 585930 338174
rect 585310 337854 585930 337938
rect 585310 337618 585342 337854
rect 585578 337618 585662 337854
rect 585898 337618 585930 337854
rect 585310 328174 585930 337618
rect 585310 327938 585342 328174
rect 585578 327938 585662 328174
rect 585898 327938 585930 328174
rect 585310 327854 585930 327938
rect 585310 327618 585342 327854
rect 585578 327618 585662 327854
rect 585898 327618 585930 327854
rect 585310 318174 585930 327618
rect 585310 317938 585342 318174
rect 585578 317938 585662 318174
rect 585898 317938 585930 318174
rect 585310 317854 585930 317938
rect 585310 317618 585342 317854
rect 585578 317618 585662 317854
rect 585898 317618 585930 317854
rect 585310 308174 585930 317618
rect 585310 307938 585342 308174
rect 585578 307938 585662 308174
rect 585898 307938 585930 308174
rect 585310 307854 585930 307938
rect 585310 307618 585342 307854
rect 585578 307618 585662 307854
rect 585898 307618 585930 307854
rect 580211 298756 580277 298757
rect 580211 298692 580212 298756
rect 580276 298692 580277 298756
rect 580211 298691 580277 298692
rect 578923 245580 578989 245581
rect 578923 245516 578924 245580
rect 578988 245516 578989 245580
rect 578923 245515 578989 245516
rect 578739 90404 578805 90405
rect 578739 90340 578740 90404
rect 578804 90340 578805 90404
rect 578739 90339 578805 90340
rect 577635 86188 577701 86189
rect 577635 86124 577636 86188
rect 577700 86124 577701 86188
rect 577635 86123 577701 86124
rect 577451 75172 577517 75173
rect 577451 75108 577452 75172
rect 577516 75108 577517 75172
rect 577451 75107 577517 75108
rect 576163 72452 576229 72453
rect 576163 72388 576164 72452
rect 576228 72388 576229 72452
rect 576163 72387 576229 72388
rect 574875 69596 574941 69597
rect 574875 69532 574876 69596
rect 574940 69532 574941 69596
rect 574875 69531 574941 69532
rect 313227 66876 313293 66877
rect 313227 66812 313228 66876
rect 313292 66812 313293 66876
rect 313227 66811 313293 66812
rect 578926 21997 578986 245515
rect 580214 89045 580274 298691
rect 585310 298174 585930 307618
rect 585310 297938 585342 298174
rect 585578 297938 585662 298174
rect 585898 297938 585930 298174
rect 585310 297854 585930 297938
rect 585310 297618 585342 297854
rect 585578 297618 585662 297854
rect 585898 297618 585930 297854
rect 585310 288174 585930 297618
rect 585310 287938 585342 288174
rect 585578 287938 585662 288174
rect 585898 287938 585930 288174
rect 585310 287854 585930 287938
rect 585310 287618 585342 287854
rect 585578 287618 585662 287854
rect 585898 287618 585930 287854
rect 585310 278174 585930 287618
rect 585310 277938 585342 278174
rect 585578 277938 585662 278174
rect 585898 277938 585930 278174
rect 585310 277854 585930 277938
rect 585310 277618 585342 277854
rect 585578 277618 585662 277854
rect 585898 277618 585930 277854
rect 585310 268174 585930 277618
rect 585310 267938 585342 268174
rect 585578 267938 585662 268174
rect 585898 267938 585930 268174
rect 585310 267854 585930 267938
rect 585310 267618 585342 267854
rect 585578 267618 585662 267854
rect 585898 267618 585930 267854
rect 580579 259452 580645 259453
rect 580579 259388 580580 259452
rect 580644 259388 580645 259452
rect 580579 259387 580645 259388
rect 580582 258909 580642 259387
rect 580579 258908 580645 258909
rect 580579 258844 580580 258908
rect 580644 258844 580645 258908
rect 580579 258843 580645 258844
rect 580582 152693 580642 258843
rect 585310 258174 585930 267618
rect 585310 257938 585342 258174
rect 585578 257938 585662 258174
rect 585898 257938 585930 258174
rect 585310 257854 585930 257938
rect 585310 257618 585342 257854
rect 585578 257618 585662 257854
rect 585898 257618 585930 257854
rect 585310 248174 585930 257618
rect 585310 247938 585342 248174
rect 585578 247938 585662 248174
rect 585898 247938 585930 248174
rect 585310 247854 585930 247938
rect 585310 247618 585342 247854
rect 585578 247618 585662 247854
rect 585898 247618 585930 247854
rect 585310 238174 585930 247618
rect 585310 237938 585342 238174
rect 585578 237938 585662 238174
rect 585898 237938 585930 238174
rect 585310 237854 585930 237938
rect 585310 237618 585342 237854
rect 585578 237618 585662 237854
rect 585898 237618 585930 237854
rect 585310 228174 585930 237618
rect 585310 227938 585342 228174
rect 585578 227938 585662 228174
rect 585898 227938 585930 228174
rect 585310 227854 585930 227938
rect 585310 227618 585342 227854
rect 585578 227618 585662 227854
rect 585898 227618 585930 227854
rect 580763 219060 580829 219061
rect 580763 218996 580764 219060
rect 580828 218996 580829 219060
rect 580763 218995 580829 218996
rect 580579 152692 580645 152693
rect 580579 152628 580580 152692
rect 580644 152628 580645 152692
rect 580579 152627 580645 152628
rect 580582 139365 580642 152627
rect 580579 139364 580645 139365
rect 580579 139300 580580 139364
rect 580644 139300 580645 139364
rect 580579 139299 580645 139300
rect 580582 112845 580642 139299
rect 580579 112844 580645 112845
rect 580579 112780 580580 112844
rect 580644 112780 580645 112844
rect 580579 112779 580645 112780
rect 580582 99517 580642 112779
rect 580579 99516 580645 99517
rect 580579 99452 580580 99516
rect 580644 99452 580645 99516
rect 580579 99451 580645 99452
rect 580211 89044 580277 89045
rect 580211 88980 580212 89044
rect 580276 88980 580277 89044
rect 580211 88979 580277 88980
rect 580582 72997 580642 99451
rect 580579 72996 580645 72997
rect 580579 72932 580580 72996
rect 580644 72932 580645 72996
rect 580579 72931 580645 72932
rect 580582 59669 580642 72931
rect 580579 59668 580645 59669
rect 580579 59604 580580 59668
rect 580644 59604 580645 59668
rect 580579 59603 580645 59604
rect 580582 33149 580642 59603
rect 580579 33148 580645 33149
rect 580579 33084 580580 33148
rect 580644 33084 580645 33148
rect 580579 33083 580645 33084
rect 578923 21996 578989 21997
rect 578923 21932 578924 21996
rect 578988 21932 578989 21996
rect 578923 21931 578989 21932
rect 306603 20636 306669 20637
rect 306603 20572 306604 20636
rect 306668 20572 306669 20636
rect 306603 20571 306669 20572
rect 311019 20636 311085 20637
rect 311019 20572 311020 20636
rect 311084 20572 311085 20636
rect 311019 20571 311085 20572
rect 580582 20501 580642 33083
rect 580579 20500 580645 20501
rect 580579 20436 580580 20500
rect 580644 20436 580645 20500
rect 580579 20435 580645 20436
rect 279003 19548 279069 19549
rect 279003 19484 279004 19548
rect 279068 19484 279069 19548
rect 279003 19483 279069 19484
rect 278635 19276 278701 19277
rect 278635 19212 278636 19276
rect 278700 19212 278701 19276
rect 278635 19211 278701 19212
rect 5027 19004 5093 19005
rect 5027 18940 5028 19004
rect 5092 18940 5093 19004
rect 5027 18939 5093 18940
rect 276427 19004 276493 19005
rect 276427 18940 276428 19004
rect 276492 18940 276493 19004
rect 276427 18939 276493 18940
rect 580766 3501 580826 218995
rect 585310 218174 585930 227618
rect 585310 217938 585342 218174
rect 585578 217938 585662 218174
rect 585898 217938 585930 218174
rect 585310 217854 585930 217938
rect 585310 217618 585342 217854
rect 585578 217618 585662 217854
rect 585898 217618 585930 217854
rect 585310 208174 585930 217618
rect 585310 207938 585342 208174
rect 585578 207938 585662 208174
rect 585898 207938 585930 208174
rect 585310 207854 585930 207938
rect 585310 207618 585342 207854
rect 585578 207618 585662 207854
rect 585898 207618 585930 207854
rect 585310 198174 585930 207618
rect 585310 197938 585342 198174
rect 585578 197938 585662 198174
rect 585898 197938 585930 198174
rect 585310 197854 585930 197938
rect 585310 197618 585342 197854
rect 585578 197618 585662 197854
rect 585898 197618 585930 197854
rect 585310 188174 585930 197618
rect 585310 187938 585342 188174
rect 585578 187938 585662 188174
rect 585898 187938 585930 188174
rect 585310 187854 585930 187938
rect 585310 187618 585342 187854
rect 585578 187618 585662 187854
rect 585898 187618 585930 187854
rect 585310 178174 585930 187618
rect 585310 177938 585342 178174
rect 585578 177938 585662 178174
rect 585898 177938 585930 178174
rect 585310 177854 585930 177938
rect 585310 177618 585342 177854
rect 585578 177618 585662 177854
rect 585898 177618 585930 177854
rect 585310 168174 585930 177618
rect 585310 167938 585342 168174
rect 585578 167938 585662 168174
rect 585898 167938 585930 168174
rect 585310 167854 585930 167938
rect 585310 167618 585342 167854
rect 585578 167618 585662 167854
rect 585898 167618 585930 167854
rect 585310 158174 585930 167618
rect 585310 157938 585342 158174
rect 585578 157938 585662 158174
rect 585898 157938 585930 158174
rect 585310 157854 585930 157938
rect 585310 157618 585342 157854
rect 585578 157618 585662 157854
rect 585898 157618 585930 157854
rect 585310 148174 585930 157618
rect 585310 147938 585342 148174
rect 585578 147938 585662 148174
rect 585898 147938 585930 148174
rect 585310 147854 585930 147938
rect 585310 147618 585342 147854
rect 585578 147618 585662 147854
rect 585898 147618 585930 147854
rect 585310 138174 585930 147618
rect 585310 137938 585342 138174
rect 585578 137938 585662 138174
rect 585898 137938 585930 138174
rect 585310 137854 585930 137938
rect 585310 137618 585342 137854
rect 585578 137618 585662 137854
rect 585898 137618 585930 137854
rect 585310 128174 585930 137618
rect 585310 127938 585342 128174
rect 585578 127938 585662 128174
rect 585898 127938 585930 128174
rect 585310 127854 585930 127938
rect 585310 127618 585342 127854
rect 585578 127618 585662 127854
rect 585898 127618 585930 127854
rect 585310 118174 585930 127618
rect 585310 117938 585342 118174
rect 585578 117938 585662 118174
rect 585898 117938 585930 118174
rect 585310 117854 585930 117938
rect 585310 117618 585342 117854
rect 585578 117618 585662 117854
rect 585898 117618 585930 117854
rect 585310 108174 585930 117618
rect 585310 107938 585342 108174
rect 585578 107938 585662 108174
rect 585898 107938 585930 108174
rect 585310 107854 585930 107938
rect 585310 107618 585342 107854
rect 585578 107618 585662 107854
rect 585898 107618 585930 107854
rect 585310 98174 585930 107618
rect 585310 97938 585342 98174
rect 585578 97938 585662 98174
rect 585898 97938 585930 98174
rect 585310 97854 585930 97938
rect 585310 97618 585342 97854
rect 585578 97618 585662 97854
rect 585898 97618 585930 97854
rect 585310 88174 585930 97618
rect 585310 87938 585342 88174
rect 585578 87938 585662 88174
rect 585898 87938 585930 88174
rect 585310 87854 585930 87938
rect 585310 87618 585342 87854
rect 585578 87618 585662 87854
rect 585898 87618 585930 87854
rect 585310 78174 585930 87618
rect 585310 77938 585342 78174
rect 585578 77938 585662 78174
rect 585898 77938 585930 78174
rect 585310 77854 585930 77938
rect 585310 77618 585342 77854
rect 585578 77618 585662 77854
rect 585898 77618 585930 77854
rect 585310 68174 585930 77618
rect 585310 67938 585342 68174
rect 585578 67938 585662 68174
rect 585898 67938 585930 68174
rect 585310 67854 585930 67938
rect 585310 67618 585342 67854
rect 585578 67618 585662 67854
rect 585898 67618 585930 67854
rect 585310 58174 585930 67618
rect 585310 57938 585342 58174
rect 585578 57938 585662 58174
rect 585898 57938 585930 58174
rect 585310 57854 585930 57938
rect 585310 57618 585342 57854
rect 585578 57618 585662 57854
rect 585898 57618 585930 57854
rect 585310 48174 585930 57618
rect 585310 47938 585342 48174
rect 585578 47938 585662 48174
rect 585898 47938 585930 48174
rect 585310 47854 585930 47938
rect 585310 47618 585342 47854
rect 585578 47618 585662 47854
rect 585898 47618 585930 47854
rect 585310 38174 585930 47618
rect 585310 37938 585342 38174
rect 585578 37938 585662 38174
rect 585898 37938 585930 38174
rect 585310 37854 585930 37938
rect 585310 37618 585342 37854
rect 585578 37618 585662 37854
rect 585898 37618 585930 37854
rect 580763 3500 580829 3501
rect 580763 3436 580764 3500
rect 580828 3436 580829 3500
rect 580763 3435 580829 3436
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 585310 -346 585930 37618
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 694454 586890 705242
rect 586270 694218 586302 694454
rect 586538 694218 586622 694454
rect 586858 694218 586890 694454
rect 586270 694134 586890 694218
rect 586270 693898 586302 694134
rect 586538 693898 586622 694134
rect 586858 693898 586890 694134
rect 586270 684454 586890 693898
rect 586270 684218 586302 684454
rect 586538 684218 586622 684454
rect 586858 684218 586890 684454
rect 586270 684134 586890 684218
rect 586270 683898 586302 684134
rect 586538 683898 586622 684134
rect 586858 683898 586890 684134
rect 586270 674454 586890 683898
rect 586270 674218 586302 674454
rect 586538 674218 586622 674454
rect 586858 674218 586890 674454
rect 586270 674134 586890 674218
rect 586270 673898 586302 674134
rect 586538 673898 586622 674134
rect 586858 673898 586890 674134
rect 586270 664454 586890 673898
rect 586270 664218 586302 664454
rect 586538 664218 586622 664454
rect 586858 664218 586890 664454
rect 586270 664134 586890 664218
rect 586270 663898 586302 664134
rect 586538 663898 586622 664134
rect 586858 663898 586890 664134
rect 586270 654454 586890 663898
rect 586270 654218 586302 654454
rect 586538 654218 586622 654454
rect 586858 654218 586890 654454
rect 586270 654134 586890 654218
rect 586270 653898 586302 654134
rect 586538 653898 586622 654134
rect 586858 653898 586890 654134
rect 586270 644454 586890 653898
rect 586270 644218 586302 644454
rect 586538 644218 586622 644454
rect 586858 644218 586890 644454
rect 586270 644134 586890 644218
rect 586270 643898 586302 644134
rect 586538 643898 586622 644134
rect 586858 643898 586890 644134
rect 586270 634454 586890 643898
rect 586270 634218 586302 634454
rect 586538 634218 586622 634454
rect 586858 634218 586890 634454
rect 586270 634134 586890 634218
rect 586270 633898 586302 634134
rect 586538 633898 586622 634134
rect 586858 633898 586890 634134
rect 586270 624454 586890 633898
rect 586270 624218 586302 624454
rect 586538 624218 586622 624454
rect 586858 624218 586890 624454
rect 586270 624134 586890 624218
rect 586270 623898 586302 624134
rect 586538 623898 586622 624134
rect 586858 623898 586890 624134
rect 586270 614454 586890 623898
rect 586270 614218 586302 614454
rect 586538 614218 586622 614454
rect 586858 614218 586890 614454
rect 586270 614134 586890 614218
rect 586270 613898 586302 614134
rect 586538 613898 586622 614134
rect 586858 613898 586890 614134
rect 586270 604454 586890 613898
rect 586270 604218 586302 604454
rect 586538 604218 586622 604454
rect 586858 604218 586890 604454
rect 586270 604134 586890 604218
rect 586270 603898 586302 604134
rect 586538 603898 586622 604134
rect 586858 603898 586890 604134
rect 586270 594454 586890 603898
rect 586270 594218 586302 594454
rect 586538 594218 586622 594454
rect 586858 594218 586890 594454
rect 586270 594134 586890 594218
rect 586270 593898 586302 594134
rect 586538 593898 586622 594134
rect 586858 593898 586890 594134
rect 586270 584454 586890 593898
rect 586270 584218 586302 584454
rect 586538 584218 586622 584454
rect 586858 584218 586890 584454
rect 586270 584134 586890 584218
rect 586270 583898 586302 584134
rect 586538 583898 586622 584134
rect 586858 583898 586890 584134
rect 586270 574454 586890 583898
rect 586270 574218 586302 574454
rect 586538 574218 586622 574454
rect 586858 574218 586890 574454
rect 586270 574134 586890 574218
rect 586270 573898 586302 574134
rect 586538 573898 586622 574134
rect 586858 573898 586890 574134
rect 586270 564454 586890 573898
rect 586270 564218 586302 564454
rect 586538 564218 586622 564454
rect 586858 564218 586890 564454
rect 586270 564134 586890 564218
rect 586270 563898 586302 564134
rect 586538 563898 586622 564134
rect 586858 563898 586890 564134
rect 586270 554454 586890 563898
rect 586270 554218 586302 554454
rect 586538 554218 586622 554454
rect 586858 554218 586890 554454
rect 586270 554134 586890 554218
rect 586270 553898 586302 554134
rect 586538 553898 586622 554134
rect 586858 553898 586890 554134
rect 586270 544454 586890 553898
rect 586270 544218 586302 544454
rect 586538 544218 586622 544454
rect 586858 544218 586890 544454
rect 586270 544134 586890 544218
rect 586270 543898 586302 544134
rect 586538 543898 586622 544134
rect 586858 543898 586890 544134
rect 586270 534454 586890 543898
rect 586270 534218 586302 534454
rect 586538 534218 586622 534454
rect 586858 534218 586890 534454
rect 586270 534134 586890 534218
rect 586270 533898 586302 534134
rect 586538 533898 586622 534134
rect 586858 533898 586890 534134
rect 586270 524454 586890 533898
rect 586270 524218 586302 524454
rect 586538 524218 586622 524454
rect 586858 524218 586890 524454
rect 586270 524134 586890 524218
rect 586270 523898 586302 524134
rect 586538 523898 586622 524134
rect 586858 523898 586890 524134
rect 586270 514454 586890 523898
rect 586270 514218 586302 514454
rect 586538 514218 586622 514454
rect 586858 514218 586890 514454
rect 586270 514134 586890 514218
rect 586270 513898 586302 514134
rect 586538 513898 586622 514134
rect 586858 513898 586890 514134
rect 586270 504454 586890 513898
rect 586270 504218 586302 504454
rect 586538 504218 586622 504454
rect 586858 504218 586890 504454
rect 586270 504134 586890 504218
rect 586270 503898 586302 504134
rect 586538 503898 586622 504134
rect 586858 503898 586890 504134
rect 586270 494454 586890 503898
rect 586270 494218 586302 494454
rect 586538 494218 586622 494454
rect 586858 494218 586890 494454
rect 586270 494134 586890 494218
rect 586270 493898 586302 494134
rect 586538 493898 586622 494134
rect 586858 493898 586890 494134
rect 586270 484454 586890 493898
rect 586270 484218 586302 484454
rect 586538 484218 586622 484454
rect 586858 484218 586890 484454
rect 586270 484134 586890 484218
rect 586270 483898 586302 484134
rect 586538 483898 586622 484134
rect 586858 483898 586890 484134
rect 586270 474454 586890 483898
rect 586270 474218 586302 474454
rect 586538 474218 586622 474454
rect 586858 474218 586890 474454
rect 586270 474134 586890 474218
rect 586270 473898 586302 474134
rect 586538 473898 586622 474134
rect 586858 473898 586890 474134
rect 586270 464454 586890 473898
rect 586270 464218 586302 464454
rect 586538 464218 586622 464454
rect 586858 464218 586890 464454
rect 586270 464134 586890 464218
rect 586270 463898 586302 464134
rect 586538 463898 586622 464134
rect 586858 463898 586890 464134
rect 586270 454454 586890 463898
rect 586270 454218 586302 454454
rect 586538 454218 586622 454454
rect 586858 454218 586890 454454
rect 586270 454134 586890 454218
rect 586270 453898 586302 454134
rect 586538 453898 586622 454134
rect 586858 453898 586890 454134
rect 586270 444454 586890 453898
rect 586270 444218 586302 444454
rect 586538 444218 586622 444454
rect 586858 444218 586890 444454
rect 586270 444134 586890 444218
rect 586270 443898 586302 444134
rect 586538 443898 586622 444134
rect 586858 443898 586890 444134
rect 586270 434454 586890 443898
rect 586270 434218 586302 434454
rect 586538 434218 586622 434454
rect 586858 434218 586890 434454
rect 586270 434134 586890 434218
rect 586270 433898 586302 434134
rect 586538 433898 586622 434134
rect 586858 433898 586890 434134
rect 586270 424454 586890 433898
rect 586270 424218 586302 424454
rect 586538 424218 586622 424454
rect 586858 424218 586890 424454
rect 586270 424134 586890 424218
rect 586270 423898 586302 424134
rect 586538 423898 586622 424134
rect 586858 423898 586890 424134
rect 586270 414454 586890 423898
rect 586270 414218 586302 414454
rect 586538 414218 586622 414454
rect 586858 414218 586890 414454
rect 586270 414134 586890 414218
rect 586270 413898 586302 414134
rect 586538 413898 586622 414134
rect 586858 413898 586890 414134
rect 586270 404454 586890 413898
rect 586270 404218 586302 404454
rect 586538 404218 586622 404454
rect 586858 404218 586890 404454
rect 586270 404134 586890 404218
rect 586270 403898 586302 404134
rect 586538 403898 586622 404134
rect 586858 403898 586890 404134
rect 586270 394454 586890 403898
rect 586270 394218 586302 394454
rect 586538 394218 586622 394454
rect 586858 394218 586890 394454
rect 586270 394134 586890 394218
rect 586270 393898 586302 394134
rect 586538 393898 586622 394134
rect 586858 393898 586890 394134
rect 586270 384454 586890 393898
rect 586270 384218 586302 384454
rect 586538 384218 586622 384454
rect 586858 384218 586890 384454
rect 586270 384134 586890 384218
rect 586270 383898 586302 384134
rect 586538 383898 586622 384134
rect 586858 383898 586890 384134
rect 586270 374454 586890 383898
rect 586270 374218 586302 374454
rect 586538 374218 586622 374454
rect 586858 374218 586890 374454
rect 586270 374134 586890 374218
rect 586270 373898 586302 374134
rect 586538 373898 586622 374134
rect 586858 373898 586890 374134
rect 586270 364454 586890 373898
rect 586270 364218 586302 364454
rect 586538 364218 586622 364454
rect 586858 364218 586890 364454
rect 586270 364134 586890 364218
rect 586270 363898 586302 364134
rect 586538 363898 586622 364134
rect 586858 363898 586890 364134
rect 586270 354454 586890 363898
rect 586270 354218 586302 354454
rect 586538 354218 586622 354454
rect 586858 354218 586890 354454
rect 586270 354134 586890 354218
rect 586270 353898 586302 354134
rect 586538 353898 586622 354134
rect 586858 353898 586890 354134
rect 586270 344454 586890 353898
rect 586270 344218 586302 344454
rect 586538 344218 586622 344454
rect 586858 344218 586890 344454
rect 586270 344134 586890 344218
rect 586270 343898 586302 344134
rect 586538 343898 586622 344134
rect 586858 343898 586890 344134
rect 586270 334454 586890 343898
rect 586270 334218 586302 334454
rect 586538 334218 586622 334454
rect 586858 334218 586890 334454
rect 586270 334134 586890 334218
rect 586270 333898 586302 334134
rect 586538 333898 586622 334134
rect 586858 333898 586890 334134
rect 586270 324454 586890 333898
rect 586270 324218 586302 324454
rect 586538 324218 586622 324454
rect 586858 324218 586890 324454
rect 586270 324134 586890 324218
rect 586270 323898 586302 324134
rect 586538 323898 586622 324134
rect 586858 323898 586890 324134
rect 586270 314454 586890 323898
rect 586270 314218 586302 314454
rect 586538 314218 586622 314454
rect 586858 314218 586890 314454
rect 586270 314134 586890 314218
rect 586270 313898 586302 314134
rect 586538 313898 586622 314134
rect 586858 313898 586890 314134
rect 586270 304454 586890 313898
rect 586270 304218 586302 304454
rect 586538 304218 586622 304454
rect 586858 304218 586890 304454
rect 586270 304134 586890 304218
rect 586270 303898 586302 304134
rect 586538 303898 586622 304134
rect 586858 303898 586890 304134
rect 586270 294454 586890 303898
rect 586270 294218 586302 294454
rect 586538 294218 586622 294454
rect 586858 294218 586890 294454
rect 586270 294134 586890 294218
rect 586270 293898 586302 294134
rect 586538 293898 586622 294134
rect 586858 293898 586890 294134
rect 586270 284454 586890 293898
rect 586270 284218 586302 284454
rect 586538 284218 586622 284454
rect 586858 284218 586890 284454
rect 586270 284134 586890 284218
rect 586270 283898 586302 284134
rect 586538 283898 586622 284134
rect 586858 283898 586890 284134
rect 586270 274454 586890 283898
rect 586270 274218 586302 274454
rect 586538 274218 586622 274454
rect 586858 274218 586890 274454
rect 586270 274134 586890 274218
rect 586270 273898 586302 274134
rect 586538 273898 586622 274134
rect 586858 273898 586890 274134
rect 586270 264454 586890 273898
rect 586270 264218 586302 264454
rect 586538 264218 586622 264454
rect 586858 264218 586890 264454
rect 586270 264134 586890 264218
rect 586270 263898 586302 264134
rect 586538 263898 586622 264134
rect 586858 263898 586890 264134
rect 586270 254454 586890 263898
rect 586270 254218 586302 254454
rect 586538 254218 586622 254454
rect 586858 254218 586890 254454
rect 586270 254134 586890 254218
rect 586270 253898 586302 254134
rect 586538 253898 586622 254134
rect 586858 253898 586890 254134
rect 586270 244454 586890 253898
rect 586270 244218 586302 244454
rect 586538 244218 586622 244454
rect 586858 244218 586890 244454
rect 586270 244134 586890 244218
rect 586270 243898 586302 244134
rect 586538 243898 586622 244134
rect 586858 243898 586890 244134
rect 586270 234454 586890 243898
rect 586270 234218 586302 234454
rect 586538 234218 586622 234454
rect 586858 234218 586890 234454
rect 586270 234134 586890 234218
rect 586270 233898 586302 234134
rect 586538 233898 586622 234134
rect 586858 233898 586890 234134
rect 586270 224454 586890 233898
rect 586270 224218 586302 224454
rect 586538 224218 586622 224454
rect 586858 224218 586890 224454
rect 586270 224134 586890 224218
rect 586270 223898 586302 224134
rect 586538 223898 586622 224134
rect 586858 223898 586890 224134
rect 586270 214454 586890 223898
rect 586270 214218 586302 214454
rect 586538 214218 586622 214454
rect 586858 214218 586890 214454
rect 586270 214134 586890 214218
rect 586270 213898 586302 214134
rect 586538 213898 586622 214134
rect 586858 213898 586890 214134
rect 586270 204454 586890 213898
rect 586270 204218 586302 204454
rect 586538 204218 586622 204454
rect 586858 204218 586890 204454
rect 586270 204134 586890 204218
rect 586270 203898 586302 204134
rect 586538 203898 586622 204134
rect 586858 203898 586890 204134
rect 586270 194454 586890 203898
rect 586270 194218 586302 194454
rect 586538 194218 586622 194454
rect 586858 194218 586890 194454
rect 586270 194134 586890 194218
rect 586270 193898 586302 194134
rect 586538 193898 586622 194134
rect 586858 193898 586890 194134
rect 586270 184454 586890 193898
rect 586270 184218 586302 184454
rect 586538 184218 586622 184454
rect 586858 184218 586890 184454
rect 586270 184134 586890 184218
rect 586270 183898 586302 184134
rect 586538 183898 586622 184134
rect 586858 183898 586890 184134
rect 586270 174454 586890 183898
rect 586270 174218 586302 174454
rect 586538 174218 586622 174454
rect 586858 174218 586890 174454
rect 586270 174134 586890 174218
rect 586270 173898 586302 174134
rect 586538 173898 586622 174134
rect 586858 173898 586890 174134
rect 586270 164454 586890 173898
rect 586270 164218 586302 164454
rect 586538 164218 586622 164454
rect 586858 164218 586890 164454
rect 586270 164134 586890 164218
rect 586270 163898 586302 164134
rect 586538 163898 586622 164134
rect 586858 163898 586890 164134
rect 586270 154454 586890 163898
rect 586270 154218 586302 154454
rect 586538 154218 586622 154454
rect 586858 154218 586890 154454
rect 586270 154134 586890 154218
rect 586270 153898 586302 154134
rect 586538 153898 586622 154134
rect 586858 153898 586890 154134
rect 586270 144454 586890 153898
rect 586270 144218 586302 144454
rect 586538 144218 586622 144454
rect 586858 144218 586890 144454
rect 586270 144134 586890 144218
rect 586270 143898 586302 144134
rect 586538 143898 586622 144134
rect 586858 143898 586890 144134
rect 586270 134454 586890 143898
rect 586270 134218 586302 134454
rect 586538 134218 586622 134454
rect 586858 134218 586890 134454
rect 586270 134134 586890 134218
rect 586270 133898 586302 134134
rect 586538 133898 586622 134134
rect 586858 133898 586890 134134
rect 586270 124454 586890 133898
rect 586270 124218 586302 124454
rect 586538 124218 586622 124454
rect 586858 124218 586890 124454
rect 586270 124134 586890 124218
rect 586270 123898 586302 124134
rect 586538 123898 586622 124134
rect 586858 123898 586890 124134
rect 586270 114454 586890 123898
rect 586270 114218 586302 114454
rect 586538 114218 586622 114454
rect 586858 114218 586890 114454
rect 586270 114134 586890 114218
rect 586270 113898 586302 114134
rect 586538 113898 586622 114134
rect 586858 113898 586890 114134
rect 586270 104454 586890 113898
rect 586270 104218 586302 104454
rect 586538 104218 586622 104454
rect 586858 104218 586890 104454
rect 586270 104134 586890 104218
rect 586270 103898 586302 104134
rect 586538 103898 586622 104134
rect 586858 103898 586890 104134
rect 586270 94454 586890 103898
rect 586270 94218 586302 94454
rect 586538 94218 586622 94454
rect 586858 94218 586890 94454
rect 586270 94134 586890 94218
rect 586270 93898 586302 94134
rect 586538 93898 586622 94134
rect 586858 93898 586890 94134
rect 586270 84454 586890 93898
rect 586270 84218 586302 84454
rect 586538 84218 586622 84454
rect 586858 84218 586890 84454
rect 586270 84134 586890 84218
rect 586270 83898 586302 84134
rect 586538 83898 586622 84134
rect 586858 83898 586890 84134
rect 586270 74454 586890 83898
rect 586270 74218 586302 74454
rect 586538 74218 586622 74454
rect 586858 74218 586890 74454
rect 586270 74134 586890 74218
rect 586270 73898 586302 74134
rect 586538 73898 586622 74134
rect 586858 73898 586890 74134
rect 586270 64454 586890 73898
rect 586270 64218 586302 64454
rect 586538 64218 586622 64454
rect 586858 64218 586890 64454
rect 586270 64134 586890 64218
rect 586270 63898 586302 64134
rect 586538 63898 586622 64134
rect 586858 63898 586890 64134
rect 586270 54454 586890 63898
rect 586270 54218 586302 54454
rect 586538 54218 586622 54454
rect 586858 54218 586890 54454
rect 586270 54134 586890 54218
rect 586270 53898 586302 54134
rect 586538 53898 586622 54134
rect 586858 53898 586890 54134
rect 586270 44454 586890 53898
rect 586270 44218 586302 44454
rect 586538 44218 586622 44454
rect 586858 44218 586890 44454
rect 586270 44134 586890 44218
rect 586270 43898 586302 44134
rect 586538 43898 586622 44134
rect 586858 43898 586890 44134
rect 586270 34454 586890 43898
rect 586270 34218 586302 34454
rect 586538 34218 586622 34454
rect 586858 34218 586890 34454
rect 586270 34134 586890 34218
rect 586270 33898 586302 34134
rect 586538 33898 586622 34134
rect 586858 33898 586890 34134
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 586270 -1306 586890 33898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 587230 -2266 587850 706202
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 588190 -3226 588810 707162
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 589150 -4186 589770 708122
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 590110 -5146 590730 709082
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 591070 -6106 591690 710042
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 592030 -7066 592650 711002
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect -2934 694218 -2698 694454
rect -2614 694218 -2378 694454
rect -2934 693898 -2698 694134
rect -2614 693898 -2378 694134
rect -2934 684218 -2698 684454
rect -2614 684218 -2378 684454
rect -2934 683898 -2698 684134
rect -2614 683898 -2378 684134
rect -2934 674218 -2698 674454
rect -2614 674218 -2378 674454
rect -2934 673898 -2698 674134
rect -2614 673898 -2378 674134
rect -2934 664218 -2698 664454
rect -2614 664218 -2378 664454
rect -2934 663898 -2698 664134
rect -2614 663898 -2378 664134
rect -2934 654218 -2698 654454
rect -2614 654218 -2378 654454
rect -2934 653898 -2698 654134
rect -2614 653898 -2378 654134
rect -2934 644218 -2698 644454
rect -2614 644218 -2378 644454
rect -2934 643898 -2698 644134
rect -2614 643898 -2378 644134
rect -2934 634218 -2698 634454
rect -2614 634218 -2378 634454
rect -2934 633898 -2698 634134
rect -2614 633898 -2378 634134
rect -2934 624218 -2698 624454
rect -2614 624218 -2378 624454
rect -2934 623898 -2698 624134
rect -2614 623898 -2378 624134
rect -2934 614218 -2698 614454
rect -2614 614218 -2378 614454
rect -2934 613898 -2698 614134
rect -2614 613898 -2378 614134
rect -2934 604218 -2698 604454
rect -2614 604218 -2378 604454
rect -2934 603898 -2698 604134
rect -2614 603898 -2378 604134
rect -2934 594218 -2698 594454
rect -2614 594218 -2378 594454
rect -2934 593898 -2698 594134
rect -2614 593898 -2378 594134
rect -2934 584218 -2698 584454
rect -2614 584218 -2378 584454
rect -2934 583898 -2698 584134
rect -2614 583898 -2378 584134
rect -2934 574218 -2698 574454
rect -2614 574218 -2378 574454
rect -2934 573898 -2698 574134
rect -2614 573898 -2378 574134
rect -2934 564218 -2698 564454
rect -2614 564218 -2378 564454
rect -2934 563898 -2698 564134
rect -2614 563898 -2378 564134
rect -2934 554218 -2698 554454
rect -2614 554218 -2378 554454
rect -2934 553898 -2698 554134
rect -2614 553898 -2378 554134
rect -2934 544218 -2698 544454
rect -2614 544218 -2378 544454
rect -2934 543898 -2698 544134
rect -2614 543898 -2378 544134
rect -2934 534218 -2698 534454
rect -2614 534218 -2378 534454
rect -2934 533898 -2698 534134
rect -2614 533898 -2378 534134
rect -2934 524218 -2698 524454
rect -2614 524218 -2378 524454
rect -2934 523898 -2698 524134
rect -2614 523898 -2378 524134
rect -2934 514218 -2698 514454
rect -2614 514218 -2378 514454
rect -2934 513898 -2698 514134
rect -2614 513898 -2378 514134
rect -2934 504218 -2698 504454
rect -2614 504218 -2378 504454
rect -2934 503898 -2698 504134
rect -2614 503898 -2378 504134
rect -2934 494218 -2698 494454
rect -2614 494218 -2378 494454
rect -2934 493898 -2698 494134
rect -2614 493898 -2378 494134
rect -2934 484218 -2698 484454
rect -2614 484218 -2378 484454
rect -2934 483898 -2698 484134
rect -2614 483898 -2378 484134
rect -2934 474218 -2698 474454
rect -2614 474218 -2378 474454
rect -2934 473898 -2698 474134
rect -2614 473898 -2378 474134
rect -2934 464218 -2698 464454
rect -2614 464218 -2378 464454
rect -2934 463898 -2698 464134
rect -2614 463898 -2378 464134
rect -2934 454218 -2698 454454
rect -2614 454218 -2378 454454
rect -2934 453898 -2698 454134
rect -2614 453898 -2378 454134
rect -2934 444218 -2698 444454
rect -2614 444218 -2378 444454
rect -2934 443898 -2698 444134
rect -2614 443898 -2378 444134
rect -2934 434218 -2698 434454
rect -2614 434218 -2378 434454
rect -2934 433898 -2698 434134
rect -2614 433898 -2378 434134
rect -2934 424218 -2698 424454
rect -2614 424218 -2378 424454
rect -2934 423898 -2698 424134
rect -2614 423898 -2378 424134
rect -2934 414218 -2698 414454
rect -2614 414218 -2378 414454
rect -2934 413898 -2698 414134
rect -2614 413898 -2378 414134
rect -2934 404218 -2698 404454
rect -2614 404218 -2378 404454
rect -2934 403898 -2698 404134
rect -2614 403898 -2378 404134
rect -2934 394218 -2698 394454
rect -2614 394218 -2378 394454
rect -2934 393898 -2698 394134
rect -2614 393898 -2378 394134
rect -2934 384218 -2698 384454
rect -2614 384218 -2378 384454
rect -2934 383898 -2698 384134
rect -2614 383898 -2378 384134
rect -2934 374218 -2698 374454
rect -2614 374218 -2378 374454
rect -2934 373898 -2698 374134
rect -2614 373898 -2378 374134
rect -2934 364218 -2698 364454
rect -2614 364218 -2378 364454
rect -2934 363898 -2698 364134
rect -2614 363898 -2378 364134
rect -2934 354218 -2698 354454
rect -2614 354218 -2378 354454
rect -2934 353898 -2698 354134
rect -2614 353898 -2378 354134
rect -2934 344218 -2698 344454
rect -2614 344218 -2378 344454
rect -2934 343898 -2698 344134
rect -2614 343898 -2378 344134
rect -2934 334218 -2698 334454
rect -2614 334218 -2378 334454
rect -2934 333898 -2698 334134
rect -2614 333898 -2378 334134
rect -2934 324218 -2698 324454
rect -2614 324218 -2378 324454
rect -2934 323898 -2698 324134
rect -2614 323898 -2378 324134
rect -2934 314218 -2698 314454
rect -2614 314218 -2378 314454
rect -2934 313898 -2698 314134
rect -2614 313898 -2378 314134
rect -2934 304218 -2698 304454
rect -2614 304218 -2378 304454
rect -2934 303898 -2698 304134
rect -2614 303898 -2378 304134
rect -2934 294218 -2698 294454
rect -2614 294218 -2378 294454
rect -2934 293898 -2698 294134
rect -2614 293898 -2378 294134
rect -2934 284218 -2698 284454
rect -2614 284218 -2378 284454
rect -2934 283898 -2698 284134
rect -2614 283898 -2378 284134
rect -2934 274218 -2698 274454
rect -2614 274218 -2378 274454
rect -2934 273898 -2698 274134
rect -2614 273898 -2378 274134
rect -2934 264218 -2698 264454
rect -2614 264218 -2378 264454
rect -2934 263898 -2698 264134
rect -2614 263898 -2378 264134
rect -2934 254218 -2698 254454
rect -2614 254218 -2378 254454
rect -2934 253898 -2698 254134
rect -2614 253898 -2378 254134
rect -2934 244218 -2698 244454
rect -2614 244218 -2378 244454
rect -2934 243898 -2698 244134
rect -2614 243898 -2378 244134
rect -2934 234218 -2698 234454
rect -2614 234218 -2378 234454
rect -2934 233898 -2698 234134
rect -2614 233898 -2378 234134
rect -2934 224218 -2698 224454
rect -2614 224218 -2378 224454
rect -2934 223898 -2698 224134
rect -2614 223898 -2378 224134
rect -2934 214218 -2698 214454
rect -2614 214218 -2378 214454
rect -2934 213898 -2698 214134
rect -2614 213898 -2378 214134
rect -2934 204218 -2698 204454
rect -2614 204218 -2378 204454
rect -2934 203898 -2698 204134
rect -2614 203898 -2378 204134
rect -2934 194218 -2698 194454
rect -2614 194218 -2378 194454
rect -2934 193898 -2698 194134
rect -2614 193898 -2378 194134
rect -2934 184218 -2698 184454
rect -2614 184218 -2378 184454
rect -2934 183898 -2698 184134
rect -2614 183898 -2378 184134
rect -2934 174218 -2698 174454
rect -2614 174218 -2378 174454
rect -2934 173898 -2698 174134
rect -2614 173898 -2378 174134
rect -2934 164218 -2698 164454
rect -2614 164218 -2378 164454
rect -2934 163898 -2698 164134
rect -2614 163898 -2378 164134
rect -2934 154218 -2698 154454
rect -2614 154218 -2378 154454
rect -2934 153898 -2698 154134
rect -2614 153898 -2378 154134
rect -2934 144218 -2698 144454
rect -2614 144218 -2378 144454
rect -2934 143898 -2698 144134
rect -2614 143898 -2378 144134
rect -2934 134218 -2698 134454
rect -2614 134218 -2378 134454
rect -2934 133898 -2698 134134
rect -2614 133898 -2378 134134
rect -2934 124218 -2698 124454
rect -2614 124218 -2378 124454
rect -2934 123898 -2698 124134
rect -2614 123898 -2378 124134
rect -2934 114218 -2698 114454
rect -2614 114218 -2378 114454
rect -2934 113898 -2698 114134
rect -2614 113898 -2378 114134
rect -2934 104218 -2698 104454
rect -2614 104218 -2378 104454
rect -2934 103898 -2698 104134
rect -2614 103898 -2378 104134
rect -2934 94218 -2698 94454
rect -2614 94218 -2378 94454
rect -2934 93898 -2698 94134
rect -2614 93898 -2378 94134
rect -2934 84218 -2698 84454
rect -2614 84218 -2378 84454
rect -2934 83898 -2698 84134
rect -2614 83898 -2378 84134
rect -2934 74218 -2698 74454
rect -2614 74218 -2378 74454
rect -2934 73898 -2698 74134
rect -2614 73898 -2378 74134
rect -2934 64218 -2698 64454
rect -2614 64218 -2378 64454
rect -2934 63898 -2698 64134
rect -2614 63898 -2378 64134
rect -2934 54218 -2698 54454
rect -2614 54218 -2378 54454
rect -2934 53898 -2698 54134
rect -2614 53898 -2378 54134
rect -2934 44218 -2698 44454
rect -2614 44218 -2378 44454
rect -2934 43898 -2698 44134
rect -2614 43898 -2378 44134
rect -2934 34218 -2698 34454
rect -2614 34218 -2378 34454
rect -2934 33898 -2698 34134
rect -2614 33898 -2378 34134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect -1974 697938 -1738 698174
rect -1654 697938 -1418 698174
rect -1974 697618 -1738 697854
rect -1654 697618 -1418 697854
rect -1974 687938 -1738 688174
rect -1654 687938 -1418 688174
rect -1974 687618 -1738 687854
rect -1654 687618 -1418 687854
rect -1974 677938 -1738 678174
rect -1654 677938 -1418 678174
rect -1974 677618 -1738 677854
rect -1654 677618 -1418 677854
rect -1974 667938 -1738 668174
rect -1654 667938 -1418 668174
rect -1974 667618 -1738 667854
rect -1654 667618 -1418 667854
rect -1974 657938 -1738 658174
rect -1654 657938 -1418 658174
rect -1974 657618 -1738 657854
rect -1654 657618 -1418 657854
rect -1974 647938 -1738 648174
rect -1654 647938 -1418 648174
rect -1974 647618 -1738 647854
rect -1654 647618 -1418 647854
rect -1974 637938 -1738 638174
rect -1654 637938 -1418 638174
rect -1974 637618 -1738 637854
rect -1654 637618 -1418 637854
rect -1974 627938 -1738 628174
rect -1654 627938 -1418 628174
rect -1974 627618 -1738 627854
rect -1654 627618 -1418 627854
rect -1974 617938 -1738 618174
rect -1654 617938 -1418 618174
rect -1974 617618 -1738 617854
rect -1654 617618 -1418 617854
rect -1974 607938 -1738 608174
rect -1654 607938 -1418 608174
rect -1974 607618 -1738 607854
rect -1654 607618 -1418 607854
rect -1974 597938 -1738 598174
rect -1654 597938 -1418 598174
rect -1974 597618 -1738 597854
rect -1654 597618 -1418 597854
rect -1974 587938 -1738 588174
rect -1654 587938 -1418 588174
rect -1974 587618 -1738 587854
rect -1654 587618 -1418 587854
rect -1974 577938 -1738 578174
rect -1654 577938 -1418 578174
rect -1974 577618 -1738 577854
rect -1654 577618 -1418 577854
rect -1974 567938 -1738 568174
rect -1654 567938 -1418 568174
rect -1974 567618 -1738 567854
rect -1654 567618 -1418 567854
rect -1974 557938 -1738 558174
rect -1654 557938 -1418 558174
rect -1974 557618 -1738 557854
rect -1654 557618 -1418 557854
rect -1974 547938 -1738 548174
rect -1654 547938 -1418 548174
rect -1974 547618 -1738 547854
rect -1654 547618 -1418 547854
rect -1974 537938 -1738 538174
rect -1654 537938 -1418 538174
rect -1974 537618 -1738 537854
rect -1654 537618 -1418 537854
rect -1974 527938 -1738 528174
rect -1654 527938 -1418 528174
rect -1974 527618 -1738 527854
rect -1654 527618 -1418 527854
rect -1974 517938 -1738 518174
rect -1654 517938 -1418 518174
rect -1974 517618 -1738 517854
rect -1654 517618 -1418 517854
rect -1974 507938 -1738 508174
rect -1654 507938 -1418 508174
rect -1974 507618 -1738 507854
rect -1654 507618 -1418 507854
rect -1974 497938 -1738 498174
rect -1654 497938 -1418 498174
rect -1974 497618 -1738 497854
rect -1654 497618 -1418 497854
rect -1974 487938 -1738 488174
rect -1654 487938 -1418 488174
rect -1974 487618 -1738 487854
rect -1654 487618 -1418 487854
rect -1974 477938 -1738 478174
rect -1654 477938 -1418 478174
rect -1974 477618 -1738 477854
rect -1654 477618 -1418 477854
rect -1974 467938 -1738 468174
rect -1654 467938 -1418 468174
rect -1974 467618 -1738 467854
rect -1654 467618 -1418 467854
rect -1974 457938 -1738 458174
rect -1654 457938 -1418 458174
rect -1974 457618 -1738 457854
rect -1654 457618 -1418 457854
rect -1974 447938 -1738 448174
rect -1654 447938 -1418 448174
rect -1974 447618 -1738 447854
rect -1654 447618 -1418 447854
rect -1974 437938 -1738 438174
rect -1654 437938 -1418 438174
rect -1974 437618 -1738 437854
rect -1654 437618 -1418 437854
rect -1974 427938 -1738 428174
rect -1654 427938 -1418 428174
rect -1974 427618 -1738 427854
rect -1654 427618 -1418 427854
rect -1974 417938 -1738 418174
rect -1654 417938 -1418 418174
rect -1974 417618 -1738 417854
rect -1654 417618 -1418 417854
rect -1974 407938 -1738 408174
rect -1654 407938 -1418 408174
rect -1974 407618 -1738 407854
rect -1654 407618 -1418 407854
rect -1974 397938 -1738 398174
rect -1654 397938 -1418 398174
rect -1974 397618 -1738 397854
rect -1654 397618 -1418 397854
rect -1974 387938 -1738 388174
rect -1654 387938 -1418 388174
rect -1974 387618 -1738 387854
rect -1654 387618 -1418 387854
rect -1974 377938 -1738 378174
rect -1654 377938 -1418 378174
rect -1974 377618 -1738 377854
rect -1654 377618 -1418 377854
rect -1974 367938 -1738 368174
rect -1654 367938 -1418 368174
rect -1974 367618 -1738 367854
rect -1654 367618 -1418 367854
rect -1974 357938 -1738 358174
rect -1654 357938 -1418 358174
rect -1974 357618 -1738 357854
rect -1654 357618 -1418 357854
rect -1974 347938 -1738 348174
rect -1654 347938 -1418 348174
rect -1974 347618 -1738 347854
rect -1654 347618 -1418 347854
rect -1974 337938 -1738 338174
rect -1654 337938 -1418 338174
rect -1974 337618 -1738 337854
rect -1654 337618 -1418 337854
rect -1974 327938 -1738 328174
rect -1654 327938 -1418 328174
rect -1974 327618 -1738 327854
rect -1654 327618 -1418 327854
rect -1974 317938 -1738 318174
rect -1654 317938 -1418 318174
rect -1974 317618 -1738 317854
rect -1654 317618 -1418 317854
rect -1974 307938 -1738 308174
rect -1654 307938 -1418 308174
rect -1974 307618 -1738 307854
rect -1654 307618 -1418 307854
rect -1974 297938 -1738 298174
rect -1654 297938 -1418 298174
rect -1974 297618 -1738 297854
rect -1654 297618 -1418 297854
rect -1974 287938 -1738 288174
rect -1654 287938 -1418 288174
rect -1974 287618 -1738 287854
rect -1654 287618 -1418 287854
rect -1974 277938 -1738 278174
rect -1654 277938 -1418 278174
rect -1974 277618 -1738 277854
rect -1654 277618 -1418 277854
rect -1974 267938 -1738 268174
rect -1654 267938 -1418 268174
rect -1974 267618 -1738 267854
rect -1654 267618 -1418 267854
rect -1974 257938 -1738 258174
rect -1654 257938 -1418 258174
rect -1974 257618 -1738 257854
rect -1654 257618 -1418 257854
rect -1974 247938 -1738 248174
rect -1654 247938 -1418 248174
rect -1974 247618 -1738 247854
rect -1654 247618 -1418 247854
rect -1974 237938 -1738 238174
rect -1654 237938 -1418 238174
rect -1974 237618 -1738 237854
rect -1654 237618 -1418 237854
rect -1974 227938 -1738 228174
rect -1654 227938 -1418 228174
rect -1974 227618 -1738 227854
rect -1654 227618 -1418 227854
rect -1974 217938 -1738 218174
rect -1654 217938 -1418 218174
rect -1974 217618 -1738 217854
rect -1654 217618 -1418 217854
rect -1974 207938 -1738 208174
rect -1654 207938 -1418 208174
rect -1974 207618 -1738 207854
rect -1654 207618 -1418 207854
rect -1974 197938 -1738 198174
rect -1654 197938 -1418 198174
rect -1974 197618 -1738 197854
rect -1654 197618 -1418 197854
rect -1974 187938 -1738 188174
rect -1654 187938 -1418 188174
rect -1974 187618 -1738 187854
rect -1654 187618 -1418 187854
rect -1974 177938 -1738 178174
rect -1654 177938 -1418 178174
rect -1974 177618 -1738 177854
rect -1654 177618 -1418 177854
rect -1974 167938 -1738 168174
rect -1654 167938 -1418 168174
rect -1974 167618 -1738 167854
rect -1654 167618 -1418 167854
rect -1974 157938 -1738 158174
rect -1654 157938 -1418 158174
rect -1974 157618 -1738 157854
rect -1654 157618 -1418 157854
rect -1974 147938 -1738 148174
rect -1654 147938 -1418 148174
rect -1974 147618 -1738 147854
rect -1654 147618 -1418 147854
rect -1974 137938 -1738 138174
rect -1654 137938 -1418 138174
rect -1974 137618 -1738 137854
rect -1654 137618 -1418 137854
rect -1974 127938 -1738 128174
rect -1654 127938 -1418 128174
rect -1974 127618 -1738 127854
rect -1654 127618 -1418 127854
rect -1974 117938 -1738 118174
rect -1654 117938 -1418 118174
rect -1974 117618 -1738 117854
rect -1654 117618 -1418 117854
rect -1974 107938 -1738 108174
rect -1654 107938 -1418 108174
rect -1974 107618 -1738 107854
rect -1654 107618 -1418 107854
rect -1974 97938 -1738 98174
rect -1654 97938 -1418 98174
rect -1974 97618 -1738 97854
rect -1654 97618 -1418 97854
rect -1974 87938 -1738 88174
rect -1654 87938 -1418 88174
rect -1974 87618 -1738 87854
rect -1654 87618 -1418 87854
rect -1974 77938 -1738 78174
rect -1654 77938 -1418 78174
rect -1974 77618 -1738 77854
rect -1654 77618 -1418 77854
rect -1974 67938 -1738 68174
rect -1654 67938 -1418 68174
rect -1974 67618 -1738 67854
rect -1654 67618 -1418 67854
rect -1974 57938 -1738 58174
rect -1654 57938 -1418 58174
rect -1974 57618 -1738 57854
rect -1654 57618 -1418 57854
rect -1974 47938 -1738 48174
rect -1654 47938 -1418 48174
rect -1974 47618 -1738 47854
rect -1654 47618 -1418 47854
rect -1974 37938 -1738 38174
rect -1654 37938 -1418 38174
rect -1974 37618 -1738 37854
rect -1654 37618 -1418 37854
rect 81714 277691 81950 277927
rect 112434 277691 112670 277927
rect 143154 277691 143390 277927
rect 149978 277691 150214 277927
rect 180698 277691 180934 277927
rect 211418 277691 211654 277927
rect 97074 274218 97310 274454
rect 97074 273898 97310 274134
rect 127794 274218 128030 274454
rect 127794 273898 128030 274134
rect 165338 274218 165574 274454
rect 165338 273898 165574 274134
rect 196058 274218 196294 274454
rect 196058 273898 196294 274134
rect 81714 267938 81950 268174
rect 81714 267618 81950 267854
rect 112434 267938 112670 268174
rect 112434 267618 112670 267854
rect 143154 267938 143390 268174
rect 143154 267618 143390 267854
rect 149978 267938 150214 268174
rect 149978 267618 150214 267854
rect 180698 267938 180934 268174
rect 180698 267618 180934 267854
rect 211418 267938 211654 268174
rect 211418 267618 211654 267854
rect 97074 264218 97310 264454
rect 97074 263898 97310 264134
rect 127794 264218 128030 264454
rect 127794 263898 128030 264134
rect 165338 264218 165574 264454
rect 165338 263898 165574 264134
rect 196058 264218 196294 264454
rect 196058 263898 196294 264134
rect 81714 257938 81950 258174
rect 81714 257618 81950 257854
rect 112434 257938 112670 258174
rect 112434 257618 112670 257854
rect 143154 257938 143390 258174
rect 143154 257618 143390 257854
rect 149978 257938 150214 258174
rect 149978 257618 150214 257854
rect 180698 257938 180934 258174
rect 180698 257618 180934 257854
rect 211418 257938 211654 258174
rect 211418 257618 211654 257854
rect 97074 254218 97310 254454
rect 97074 253898 97310 254134
rect 127794 254218 128030 254454
rect 127794 253898 128030 254134
rect 165338 254218 165574 254454
rect 165338 253898 165574 254134
rect 196058 254218 196294 254454
rect 196058 253898 196294 254134
rect 81714 247938 81950 248174
rect 81714 247618 81950 247854
rect 112434 247938 112670 248174
rect 112434 247618 112670 247854
rect 143154 247938 143390 248174
rect 143154 247618 143390 247854
rect 149978 247938 150214 248174
rect 149978 247618 150214 247854
rect 180698 247938 180934 248174
rect 180698 247618 180934 247854
rect 211418 247938 211654 248174
rect 211418 247618 211654 247854
rect 97074 244218 97310 244454
rect 97074 243898 97310 244134
rect 127794 244218 128030 244454
rect 127794 243898 128030 244134
rect 165338 244218 165574 244454
rect 165338 243898 165574 244134
rect 196058 244218 196294 244454
rect 196058 243898 196294 244134
rect 81714 237938 81950 238174
rect 81714 237618 81950 237854
rect 112434 237938 112670 238174
rect 112434 237618 112670 237854
rect 143154 237938 143390 238174
rect 143154 237618 143390 237854
rect 149978 237938 150214 238174
rect 149978 237618 150214 237854
rect 180698 237938 180934 238174
rect 180698 237618 180934 237854
rect 211418 237938 211654 238174
rect 211418 237618 211654 237854
rect 14107 207938 14343 208174
rect 14107 207618 14343 207854
rect 21949 207938 22185 208174
rect 21949 207618 22185 207854
rect 29791 207938 30027 208174
rect 29791 207618 30027 207854
rect 37633 207938 37869 208174
rect 37633 207618 37869 207854
rect 42310 207938 42546 208174
rect 42630 207938 42866 208174
rect 42950 207938 43186 208174
rect 42310 207618 42546 207854
rect 42630 207618 42866 207854
rect 42950 207618 43186 207854
rect 18028 204218 18264 204454
rect 18028 203898 18264 204134
rect 25870 204218 26106 204454
rect 25870 203898 26106 204134
rect 33712 204218 33948 204454
rect 33712 203898 33948 204134
rect 41554 204218 41790 204454
rect 41554 203898 41790 204134
rect 52160 204218 52396 204454
rect 52160 203898 52396 204134
rect 60002 204218 60238 204454
rect 60002 203898 60238 204134
rect 67844 204218 68080 204454
rect 67844 203898 68080 204134
rect 75686 204218 75922 204454
rect 75686 203898 75922 204134
rect 14107 197938 14343 198174
rect 14107 197618 14343 197854
rect 21949 197938 22185 198174
rect 21949 197618 22185 197854
rect 29791 197938 30027 198174
rect 29791 197618 30027 197854
rect 37633 197938 37869 198174
rect 37633 197618 37869 197854
rect 42310 197938 42546 198174
rect 42630 197938 42866 198174
rect 42950 197938 43186 198174
rect 42310 197618 42546 197854
rect 42630 197618 42866 197854
rect 42950 197618 43186 197854
rect 18028 194218 18264 194454
rect 18028 193898 18264 194134
rect 25870 194218 26106 194454
rect 25870 193898 26106 194134
rect 33712 194218 33948 194454
rect 33712 193898 33948 194134
rect 41554 194218 41790 194454
rect 41554 193898 41790 194134
rect 52160 194218 52396 194454
rect 52160 193898 52396 194134
rect 60002 194218 60238 194454
rect 60002 193898 60238 194134
rect 67844 194218 68080 194454
rect 67844 193898 68080 194134
rect 75686 194218 75922 194454
rect 75686 193898 75922 194134
rect 116503 227938 116739 228174
rect 116503 227618 116739 227854
rect 124345 227938 124581 228174
rect 124345 227618 124581 227854
rect 132187 227938 132423 228174
rect 132187 227618 132423 227854
rect 140029 227938 140265 228174
rect 140029 227618 140265 227854
rect 120424 224218 120660 224454
rect 120424 223898 120660 224134
rect 128266 224218 128502 224454
rect 128266 223898 128502 224134
rect 136108 224218 136344 224454
rect 136108 223898 136344 224134
rect 143950 224218 144186 224454
rect 143950 223898 144186 224134
rect 116503 217938 116739 218174
rect 116503 217618 116739 217854
rect 124345 217938 124581 218174
rect 124345 217618 124581 217854
rect 132187 217938 132423 218174
rect 132187 217618 132423 217854
rect 140029 217938 140265 218174
rect 140029 217618 140265 217854
rect 120424 214218 120660 214454
rect 120424 213898 120660 214134
rect 128266 214218 128502 214454
rect 128266 213898 128502 214134
rect 136108 214218 136344 214454
rect 136108 213898 136344 214134
rect 143950 214218 144186 214454
rect 143950 213898 144186 214134
rect 116503 207938 116739 208174
rect 116503 207618 116739 207854
rect 124345 207938 124581 208174
rect 124345 207618 124581 207854
rect 132187 207938 132423 208174
rect 132187 207618 132423 207854
rect 140029 207938 140265 208174
rect 140029 207618 140265 207854
rect 120424 204218 120660 204454
rect 120424 203898 120660 204134
rect 128266 204218 128502 204454
rect 128266 203898 128502 204134
rect 136108 204218 136344 204454
rect 136108 203898 136344 204134
rect 143950 204218 144186 204454
rect 143950 203898 144186 204134
rect 116503 197938 116739 198174
rect 116503 197618 116739 197854
rect 124345 197938 124581 198174
rect 124345 197618 124581 197854
rect 132187 197938 132423 198174
rect 132187 197618 132423 197854
rect 140029 197938 140265 198174
rect 140029 197618 140265 197854
rect 120424 194218 120660 194454
rect 120424 193898 120660 194134
rect 128266 194218 128502 194454
rect 128266 193898 128502 194134
rect 136108 194218 136344 194454
rect 136108 193898 136344 194134
rect 143950 194218 144186 194454
rect 143950 193898 144186 194134
rect 184767 207938 185003 208174
rect 184767 207618 185003 207854
rect 192609 207938 192845 208174
rect 192609 207618 192845 207854
rect 200451 207938 200687 208174
rect 200451 207618 200687 207854
rect 208293 207938 208529 208174
rect 208293 207618 208529 207854
rect 218899 207938 219135 208174
rect 218899 207618 219135 207854
rect 226741 207938 226977 208174
rect 226741 207618 226977 207854
rect 234583 207938 234819 208174
rect 234583 207618 234819 207854
rect 242425 207938 242661 208174
rect 242425 207618 242661 207854
rect 253031 207938 253267 208174
rect 253031 207618 253267 207854
rect 260873 207938 261109 208174
rect 260873 207618 261109 207854
rect 268715 207938 268951 208174
rect 268715 207618 268951 207854
rect 276557 207938 276793 208174
rect 276557 207618 276793 207854
rect 188688 204218 188924 204454
rect 188688 203898 188924 204134
rect 196530 204218 196766 204454
rect 196530 203898 196766 204134
rect 204372 204218 204608 204454
rect 204372 203898 204608 204134
rect 212214 204218 212450 204454
rect 212214 203898 212450 204134
rect 222820 204218 223056 204454
rect 222820 203898 223056 204134
rect 230662 204218 230898 204454
rect 230662 203898 230898 204134
rect 238504 204218 238740 204454
rect 238504 203898 238740 204134
rect 246346 204218 246582 204454
rect 246346 203898 246582 204134
rect 256952 204218 257188 204454
rect 256952 203898 257188 204134
rect 264794 204218 265030 204454
rect 264794 203898 265030 204134
rect 272636 204218 272872 204454
rect 272636 203898 272872 204134
rect 280478 204218 280714 204454
rect 280478 203898 280714 204134
rect 184767 197938 185003 198174
rect 184767 197618 185003 197854
rect 192609 197938 192845 198174
rect 192609 197618 192845 197854
rect 200451 197938 200687 198174
rect 200451 197618 200687 197854
rect 208293 197938 208529 198174
rect 208293 197618 208529 197854
rect 218899 197938 219135 198174
rect 218899 197618 219135 197854
rect 226741 197938 226977 198174
rect 226741 197618 226977 197854
rect 234583 197938 234819 198174
rect 234583 197618 234819 197854
rect 242425 197938 242661 198174
rect 242425 197618 242661 197854
rect 253031 197938 253267 198174
rect 253031 197618 253267 197854
rect 260873 197938 261109 198174
rect 260873 197618 261109 197854
rect 268715 197938 268951 198174
rect 268715 197618 268951 197854
rect 276557 197938 276793 198174
rect 276557 197618 276793 197854
rect 188688 194218 188924 194454
rect 188688 193898 188924 194134
rect 196530 194218 196766 194454
rect 196530 193898 196766 194134
rect 204372 194218 204608 194454
rect 204372 193898 204608 194134
rect 212214 194218 212450 194454
rect 212214 193898 212450 194134
rect 222820 194218 223056 194454
rect 222820 193898 223056 194134
rect 230662 194218 230898 194454
rect 230662 193898 230898 194134
rect 238504 194218 238740 194454
rect 238504 193898 238740 194134
rect 246346 194218 246582 194454
rect 246346 193898 246582 194134
rect 256952 194218 257188 194454
rect 256952 193898 257188 194134
rect 264794 194218 265030 194454
rect 264794 193898 265030 194134
rect 272636 194218 272872 194454
rect 272636 193898 272872 194134
rect 280478 194218 280714 194454
rect 280478 193898 280714 194134
rect 43984 187938 44220 188174
rect 43984 187618 44220 187854
rect 111581 187938 111817 188174
rect 111581 187618 111817 187854
rect 179178 187938 179414 188174
rect 179178 187618 179414 187854
rect 246775 187938 247011 188174
rect 246775 187618 247011 187854
rect 77782 184218 78018 184454
rect 77782 183898 78018 184134
rect 145379 184218 145615 184454
rect 145379 183898 145615 184134
rect 212976 184218 213212 184454
rect 212976 183898 213212 184134
rect 280573 184218 280809 184454
rect 280573 183898 280809 184134
rect 48239 177643 48475 177879
rect 56081 177643 56317 177879
rect 63923 177643 64159 177879
rect 71765 177643 72001 177879
rect 82371 177643 82607 177879
rect 90213 177643 90449 177879
rect 98055 177643 98291 177879
rect 105897 177643 106133 177879
rect 116503 177643 116739 177879
rect 124345 177643 124581 177879
rect 132187 177643 132423 177879
rect 140029 177643 140265 177879
rect 149978 177643 150214 177879
rect 180698 177643 180934 177879
rect 211418 177643 211654 177879
rect 242138 177643 242374 177879
rect 272858 177643 273094 177879
rect 52160 174218 52396 174454
rect 52160 173898 52396 174134
rect 60002 174218 60238 174454
rect 60002 173898 60238 174134
rect 67844 174218 68080 174454
rect 67844 173898 68080 174134
rect 75686 174218 75922 174454
rect 75686 173898 75922 174134
rect 86292 174218 86528 174454
rect 86292 173898 86528 174134
rect 94134 174218 94370 174454
rect 94134 173898 94370 174134
rect 101976 174218 102212 174454
rect 101976 173898 102212 174134
rect 109818 174218 110054 174454
rect 109818 173898 110054 174134
rect 120424 174218 120660 174454
rect 120424 173898 120660 174134
rect 128266 174218 128502 174454
rect 128266 173898 128502 174134
rect 136108 174218 136344 174454
rect 136108 173898 136344 174134
rect 143950 174218 144186 174454
rect 143950 173898 144186 174134
rect 165338 174218 165574 174454
rect 165338 173898 165574 174134
rect 196058 174218 196294 174454
rect 196058 173898 196294 174134
rect 226778 174218 227014 174454
rect 226778 173898 227014 174134
rect 257498 174218 257734 174454
rect 257498 173898 257734 174134
rect 48239 167938 48475 168174
rect 48239 167618 48475 167854
rect 56081 167938 56317 168174
rect 56081 167618 56317 167854
rect 63923 167938 64159 168174
rect 63923 167618 64159 167854
rect 71765 167938 72001 168174
rect 71765 167618 72001 167854
rect 82371 167938 82607 168174
rect 82371 167618 82607 167854
rect 90213 167938 90449 168174
rect 90213 167618 90449 167854
rect 98055 167938 98291 168174
rect 98055 167618 98291 167854
rect 105897 167938 106133 168174
rect 105897 167618 106133 167854
rect 116503 167938 116739 168174
rect 116503 167618 116739 167854
rect 124345 167938 124581 168174
rect 124345 167618 124581 167854
rect 132187 167938 132423 168174
rect 132187 167618 132423 167854
rect 140029 167938 140265 168174
rect 140029 167618 140265 167854
rect 149978 167938 150214 168174
rect 149978 167618 150214 167854
rect 180698 167938 180934 168174
rect 180698 167618 180934 167854
rect 211418 167938 211654 168174
rect 211418 167618 211654 167854
rect 242138 167938 242374 168174
rect 242138 167618 242374 167854
rect 272858 167938 273094 168174
rect 272858 167618 273094 167854
rect 52160 164218 52396 164454
rect 52160 163898 52396 164134
rect 60002 164218 60238 164454
rect 60002 163898 60238 164134
rect 67844 164218 68080 164454
rect 67844 163898 68080 164134
rect 75686 164218 75922 164454
rect 75686 163898 75922 164134
rect 86292 164218 86528 164454
rect 86292 163898 86528 164134
rect 94134 164218 94370 164454
rect 94134 163898 94370 164134
rect 101976 164218 102212 164454
rect 101976 163898 102212 164134
rect 109818 164218 110054 164454
rect 109818 163898 110054 164134
rect 120424 164218 120660 164454
rect 120424 163898 120660 164134
rect 128266 164218 128502 164454
rect 128266 163898 128502 164134
rect 136108 164218 136344 164454
rect 136108 163898 136344 164134
rect 143950 164218 144186 164454
rect 143950 163898 144186 164134
rect 165338 164218 165574 164454
rect 165338 163898 165574 164134
rect 196058 164218 196294 164454
rect 196058 163898 196294 164134
rect 226778 164218 227014 164454
rect 226778 163898 227014 164134
rect 257498 164218 257734 164454
rect 257498 163898 257734 164134
rect 277814 164218 278050 164454
rect 277814 163898 278050 164134
rect 48239 157938 48475 158174
rect 48239 157618 48475 157854
rect 56081 157938 56317 158174
rect 56081 157618 56317 157854
rect 63923 157938 64159 158174
rect 63923 157618 64159 157854
rect 71765 157938 72001 158174
rect 71765 157618 72001 157854
rect 82371 157938 82607 158174
rect 82371 157618 82607 157854
rect 90213 157938 90449 158174
rect 90213 157618 90449 157854
rect 98055 157938 98291 158174
rect 98055 157618 98291 157854
rect 105897 157938 106133 158174
rect 105897 157618 106133 157854
rect 149978 157938 150214 158174
rect 149978 157618 150214 157854
rect 180698 157938 180934 158174
rect 180698 157618 180934 157854
rect 277262 157938 277498 158174
rect 277262 157618 277498 157854
rect 52160 154218 52396 154454
rect 52160 153898 52396 154134
rect 60002 154218 60238 154454
rect 60002 153898 60238 154134
rect 67844 154218 68080 154454
rect 67844 153898 68080 154134
rect 75686 154218 75922 154454
rect 75686 153898 75922 154134
rect 86292 154218 86528 154454
rect 86292 153898 86528 154134
rect 94134 154218 94370 154454
rect 94134 153898 94370 154134
rect 101976 154218 102212 154454
rect 101976 153898 102212 154134
rect 109818 154218 110054 154454
rect 109818 153898 110054 154134
rect 165338 154218 165574 154454
rect 165338 153898 165574 154134
rect 277814 154218 278050 154454
rect 277814 153898 278050 154134
rect 48239 147938 48475 148174
rect 48239 147618 48475 147854
rect 56081 147938 56317 148174
rect 56081 147618 56317 147854
rect 63923 147938 64159 148174
rect 63923 147618 64159 147854
rect 71765 147938 72001 148174
rect 71765 147618 72001 147854
rect 82371 147938 82607 148174
rect 82371 147618 82607 147854
rect 90213 147938 90449 148174
rect 90213 147618 90449 147854
rect 98055 147938 98291 148174
rect 98055 147618 98291 147854
rect 105897 147938 106133 148174
rect 105897 147618 106133 147854
rect 149978 147938 150214 148174
rect 149978 147618 150214 147854
rect 180698 147938 180934 148174
rect 180698 147618 180934 147854
rect 277262 147938 277498 148174
rect 277262 147618 277498 147854
rect 52160 144218 52396 144454
rect 52160 143898 52396 144134
rect 60002 144218 60238 144454
rect 60002 143898 60238 144134
rect 67844 144218 68080 144454
rect 67844 143898 68080 144134
rect 75686 144218 75922 144454
rect 75686 143898 75922 144134
rect 86292 144218 86528 144454
rect 86292 143898 86528 144134
rect 94134 144218 94370 144454
rect 94134 143898 94370 144134
rect 101976 144218 102212 144454
rect 101976 143898 102212 144134
rect 109818 144218 110054 144454
rect 109818 143898 110054 144134
rect 165338 144218 165574 144454
rect 165338 143898 165574 144134
rect 277814 144218 278050 144454
rect 277814 143898 278050 144134
rect 48239 137938 48475 138174
rect 48239 137618 48475 137854
rect 56081 137938 56317 138174
rect 56081 137618 56317 137854
rect 63923 137938 64159 138174
rect 63923 137618 64159 137854
rect 71765 137938 72001 138174
rect 71765 137618 72001 137854
rect 82371 137938 82607 138174
rect 82371 137618 82607 137854
rect 90213 137938 90449 138174
rect 90213 137618 90449 137854
rect 98055 137938 98291 138174
rect 98055 137618 98291 137854
rect 105897 137938 106133 138174
rect 105897 137618 106133 137854
rect 149978 137938 150214 138174
rect 149978 137618 150214 137854
rect 180698 137938 180934 138174
rect 180698 137618 180934 137854
rect 211418 137938 211654 138174
rect 211418 137618 211654 137854
rect 242138 137938 242374 138174
rect 242138 137618 242374 137854
rect 272858 137938 273094 138174
rect 272858 137618 273094 137854
rect 277262 137938 277498 138174
rect 277262 137618 277498 137854
rect 13450 127938 13686 128174
rect 13450 127618 13686 127854
rect 44170 127938 44406 128174
rect 44170 127618 44406 127854
rect 74890 127938 75126 128174
rect 74890 127618 75126 127854
rect 105610 127938 105846 128174
rect 105610 127618 105846 127854
rect 136330 127938 136566 128174
rect 136330 127618 136566 127854
rect 167050 127938 167286 128174
rect 167050 127618 167286 127854
rect 197770 127938 198006 128174
rect 197770 127618 198006 127854
rect 228490 127938 228726 128174
rect 228490 127618 228726 127854
rect 259210 127938 259446 128174
rect 259210 127618 259446 127854
rect 28810 124218 29046 124454
rect 28810 123898 29046 124134
rect 59530 124218 59766 124454
rect 59530 123898 59766 124134
rect 90250 124218 90486 124454
rect 90250 123898 90486 124134
rect 120970 124218 121206 124454
rect 120970 123898 121206 124134
rect 151690 124218 151926 124454
rect 151690 123898 151926 124134
rect 182410 124218 182646 124454
rect 182410 123898 182646 124134
rect 213130 124218 213366 124454
rect 213130 123898 213366 124134
rect 243850 124218 244086 124454
rect 243850 123898 244086 124134
rect 274570 124218 274806 124454
rect 274570 123898 274806 124134
rect 13450 117938 13686 118174
rect 13450 117618 13686 117854
rect 44170 117938 44406 118174
rect 44170 117618 44406 117854
rect 74890 117938 75126 118174
rect 74890 117618 75126 117854
rect 105610 117938 105846 118174
rect 105610 117618 105846 117854
rect 136330 117938 136566 118174
rect 136330 117618 136566 117854
rect 167050 117938 167286 118174
rect 167050 117618 167286 117854
rect 197770 117938 198006 118174
rect 197770 117618 198006 117854
rect 228490 117938 228726 118174
rect 228490 117618 228726 117854
rect 259210 117938 259446 118174
rect 259210 117618 259446 117854
rect 28810 114218 29046 114454
rect 28810 113898 29046 114134
rect 59530 114218 59766 114454
rect 59530 113898 59766 114134
rect 90250 114218 90486 114454
rect 90250 113898 90486 114134
rect 120970 114218 121206 114454
rect 120970 113898 121206 114134
rect 151690 114218 151926 114454
rect 151690 113898 151926 114134
rect 182410 114218 182646 114454
rect 182410 113898 182646 114134
rect 213130 114218 213366 114454
rect 213130 113898 213366 114134
rect 243850 114218 244086 114454
rect 243850 113898 244086 114134
rect 274570 114218 274806 114454
rect 274570 113898 274806 114134
rect 13450 107938 13686 108174
rect 13450 107618 13686 107854
rect 44170 107938 44406 108174
rect 44170 107618 44406 107854
rect 74890 107938 75126 108174
rect 74890 107618 75126 107854
rect 105610 107938 105846 108174
rect 105610 107618 105846 107854
rect 136330 107938 136566 108174
rect 136330 107618 136566 107854
rect 167050 107938 167286 108174
rect 167050 107618 167286 107854
rect 197770 107938 198006 108174
rect 197770 107618 198006 107854
rect 228490 107938 228726 108174
rect 228490 107618 228726 107854
rect 259210 107938 259446 108174
rect 259210 107618 259446 107854
rect 28810 104218 29046 104454
rect 28810 103898 29046 104134
rect 59530 104218 59766 104454
rect 59530 103898 59766 104134
rect 90250 104218 90486 104454
rect 90250 103898 90486 104134
rect 120970 104218 121206 104454
rect 120970 103898 121206 104134
rect 151690 104218 151926 104454
rect 151690 103898 151926 104134
rect 182410 104218 182646 104454
rect 182410 103898 182646 104134
rect 213130 104218 213366 104454
rect 213130 103898 213366 104134
rect 243850 104218 244086 104454
rect 243850 103898 244086 104134
rect 274570 104218 274806 104454
rect 274570 103898 274806 104134
rect 13450 97938 13686 98174
rect 13450 97618 13686 97854
rect 44170 97938 44406 98174
rect 44170 97618 44406 97854
rect 74890 97938 75126 98174
rect 74890 97618 75126 97854
rect 105610 97938 105846 98174
rect 105610 97618 105846 97854
rect 136330 97938 136566 98174
rect 136330 97618 136566 97854
rect 167050 97938 167286 98174
rect 167050 97618 167286 97854
rect 197770 97938 198006 98174
rect 197770 97618 198006 97854
rect 228490 97938 228726 98174
rect 228490 97618 228726 97854
rect 259210 97938 259446 98174
rect 259210 97618 259446 97854
rect 28810 94218 29046 94454
rect 28810 93898 29046 94134
rect 59530 94218 59766 94454
rect 59530 93898 59766 94134
rect 90250 94218 90486 94454
rect 90250 93898 90486 94134
rect 120970 94218 121206 94454
rect 120970 93898 121206 94134
rect 151690 94218 151926 94454
rect 151690 93898 151926 94134
rect 182410 94218 182646 94454
rect 182410 93898 182646 94134
rect 213130 94218 213366 94454
rect 213130 93898 213366 94134
rect 243850 94218 244086 94454
rect 243850 93898 244086 94134
rect 274570 94218 274806 94454
rect 274570 93898 274806 94134
rect 585342 697938 585578 698174
rect 585662 697938 585898 698174
rect 585342 697618 585578 697854
rect 585662 697618 585898 697854
rect 585342 687938 585578 688174
rect 585662 687938 585898 688174
rect 585342 687618 585578 687854
rect 585662 687618 585898 687854
rect 585342 677938 585578 678174
rect 585662 677938 585898 678174
rect 585342 677618 585578 677854
rect 585662 677618 585898 677854
rect 303504 317938 303740 318174
rect 303504 317618 303740 317854
rect 437872 317938 438108 318174
rect 437872 317618 438108 317854
rect 302824 314218 303060 314454
rect 302824 313898 303060 314134
rect 438552 314218 438788 314454
rect 438552 313898 438788 314134
rect 303504 307938 303740 308174
rect 303504 307618 303740 307854
rect 437872 307938 438108 308174
rect 437872 307618 438108 307854
rect 302824 304218 303060 304454
rect 302824 303898 303060 304134
rect 438552 304218 438788 304454
rect 438552 303898 438788 304134
rect 303504 297938 303740 298174
rect 303504 297618 303740 297854
rect 437872 297938 438108 298174
rect 437872 297618 438108 297854
rect 302824 294218 303060 294454
rect 302824 293898 303060 294134
rect 438552 294218 438788 294454
rect 438552 293898 438788 294134
rect 303504 287938 303740 288174
rect 303504 287618 303740 287854
rect 437872 287938 438108 288174
rect 437872 287618 438108 287854
rect 302824 284218 303060 284454
rect 302824 283898 303060 284134
rect 438552 284218 438788 284454
rect 438552 283898 438788 284134
rect 303504 277938 303740 278174
rect 303504 277618 303740 277854
rect 437872 277938 438108 278174
rect 437872 277618 438108 277854
rect 302824 274218 303060 274454
rect 302824 273898 303060 274134
rect 438552 274218 438788 274454
rect 438552 273898 438788 274134
rect 303504 267938 303740 268174
rect 303504 267618 303740 267854
rect 437872 267938 438108 268174
rect 437872 267618 438108 267854
rect 302824 264218 303060 264454
rect 302824 263898 303060 264134
rect 438552 264218 438788 264454
rect 438552 263898 438788 264134
rect 303504 257938 303740 258174
rect 303504 257618 303740 257854
rect 437872 257938 438108 258174
rect 437872 257618 438108 257854
rect 302824 254218 303060 254454
rect 302824 253898 303060 254134
rect 438552 254218 438788 254454
rect 438552 253898 438788 254134
rect 303504 247938 303740 248174
rect 303504 247618 303740 247854
rect 437872 247938 438108 248174
rect 437872 247618 438108 247854
rect 302824 244218 303060 244454
rect 302824 243898 303060 244134
rect 438552 244218 438788 244454
rect 438552 243898 438788 244134
rect 307407 207938 307643 208174
rect 307407 207618 307643 207854
rect 315249 207938 315485 208174
rect 315249 207618 315485 207854
rect 323091 207938 323327 208174
rect 323091 207618 323327 207854
rect 330933 207938 331169 208174
rect 330933 207618 331169 207854
rect 303486 204218 303722 204454
rect 303486 203898 303722 204134
rect 311328 204218 311564 204454
rect 311328 203898 311564 204134
rect 319170 204218 319406 204454
rect 319170 203898 319406 204134
rect 327012 204218 327248 204454
rect 327012 203898 327248 204134
rect 307407 197938 307643 198174
rect 307407 197618 307643 197854
rect 315249 197938 315485 198174
rect 315249 197618 315485 197854
rect 323091 197938 323327 198174
rect 323091 197618 323327 197854
rect 330933 197938 331169 198174
rect 330933 197618 331169 197854
rect 303486 194218 303722 194454
rect 303486 193898 303722 194134
rect 311328 194218 311564 194454
rect 311328 193898 311564 194134
rect 319170 194218 319406 194454
rect 319170 193898 319406 194134
rect 327012 194218 327248 194454
rect 327012 193898 327248 194134
rect 409803 227938 410039 228174
rect 409803 227618 410039 227854
rect 417645 227938 417881 228174
rect 417645 227618 417881 227854
rect 425487 227938 425723 228174
rect 425487 227618 425723 227854
rect 433329 227938 433565 228174
rect 433329 227618 433565 227854
rect 405882 224218 406118 224454
rect 405882 223898 406118 224134
rect 413724 224218 413960 224454
rect 413724 223898 413960 224134
rect 421566 224218 421802 224454
rect 421566 223898 421802 224134
rect 429408 224218 429644 224454
rect 429408 223898 429644 224134
rect 409803 217938 410039 218174
rect 409803 217618 410039 217854
rect 417645 217938 417881 218174
rect 417645 217618 417881 217854
rect 425487 217938 425723 218174
rect 425487 217618 425723 217854
rect 433329 217938 433565 218174
rect 433329 217618 433565 217854
rect 405882 214218 406118 214454
rect 405882 213898 406118 214134
rect 413724 214218 413960 214454
rect 413724 213898 413960 214134
rect 421566 214218 421802 214454
rect 421566 213898 421802 214134
rect 429408 214218 429644 214454
rect 429408 213898 429644 214134
rect 341539 207938 341775 208174
rect 341539 207618 341775 207854
rect 349381 207938 349617 208174
rect 349381 207618 349617 207854
rect 357223 207938 357459 208174
rect 357223 207618 357459 207854
rect 365065 207938 365301 208174
rect 365065 207618 365301 207854
rect 375671 207938 375907 208174
rect 375671 207618 375907 207854
rect 383513 207938 383749 208174
rect 383513 207618 383749 207854
rect 391355 207938 391591 208174
rect 391355 207618 391591 207854
rect 399197 207938 399433 208174
rect 399197 207618 399433 207854
rect 409803 207938 410039 208174
rect 409803 207618 410039 207854
rect 417645 207938 417881 208174
rect 417645 207618 417881 207854
rect 425487 207938 425723 208174
rect 425487 207618 425723 207854
rect 433329 207938 433565 208174
rect 433329 207618 433565 207854
rect 443935 207938 444171 208174
rect 443935 207618 444171 207854
rect 451777 207938 452013 208174
rect 451777 207618 452013 207854
rect 459619 207938 459855 208174
rect 459619 207618 459855 207854
rect 467461 207938 467697 208174
rect 467461 207618 467697 207854
rect 478067 207938 478303 208174
rect 478067 207618 478303 207854
rect 485909 207938 486145 208174
rect 485909 207618 486145 207854
rect 493751 207938 493987 208174
rect 493751 207618 493987 207854
rect 501593 207938 501829 208174
rect 501593 207618 501829 207854
rect 512199 207938 512435 208174
rect 512199 207618 512435 207854
rect 520041 207938 520277 208174
rect 520041 207618 520277 207854
rect 527883 207938 528119 208174
rect 527883 207618 528119 207854
rect 535725 207938 535961 208174
rect 535725 207618 535961 207854
rect 546331 207938 546567 208174
rect 546331 207618 546567 207854
rect 554173 207938 554409 208174
rect 554173 207618 554409 207854
rect 562015 207938 562251 208174
rect 562015 207618 562251 207854
rect 569857 207938 570093 208174
rect 569857 207618 570093 207854
rect 337618 204218 337854 204454
rect 337618 203898 337854 204134
rect 345460 204218 345696 204454
rect 345460 203898 345696 204134
rect 353302 204218 353538 204454
rect 353302 203898 353538 204134
rect 361144 204218 361380 204454
rect 361144 203898 361380 204134
rect 371750 204218 371986 204454
rect 371750 203898 371986 204134
rect 379592 204218 379828 204454
rect 379592 203898 379828 204134
rect 387434 204218 387670 204454
rect 387434 203898 387670 204134
rect 395276 204218 395512 204454
rect 395276 203898 395512 204134
rect 405882 204218 406118 204454
rect 405882 203898 406118 204134
rect 413724 204218 413960 204454
rect 413724 203898 413960 204134
rect 421566 204218 421802 204454
rect 421566 203898 421802 204134
rect 429408 204218 429644 204454
rect 429408 203898 429644 204134
rect 440014 204218 440250 204454
rect 440014 203898 440250 204134
rect 447856 204218 448092 204454
rect 447856 203898 448092 204134
rect 455698 204218 455934 204454
rect 455698 203898 455934 204134
rect 463540 204218 463776 204454
rect 463540 203898 463776 204134
rect 474146 204218 474382 204454
rect 474146 203898 474382 204134
rect 481988 204218 482224 204454
rect 481988 203898 482224 204134
rect 489830 204218 490066 204454
rect 489830 203898 490066 204134
rect 497672 204218 497908 204454
rect 497672 203898 497908 204134
rect 508278 204218 508514 204454
rect 508278 203898 508514 204134
rect 516120 204218 516356 204454
rect 516120 203898 516356 204134
rect 523962 204218 524198 204454
rect 523962 203898 524198 204134
rect 531804 204218 532040 204454
rect 531804 203898 532040 204134
rect 542410 204218 542646 204454
rect 542410 203898 542646 204134
rect 550252 204218 550488 204454
rect 550252 203898 550488 204134
rect 558094 204218 558330 204454
rect 558094 203898 558330 204134
rect 565936 204218 566172 204454
rect 565936 203898 566172 204134
rect 341539 197938 341775 198174
rect 341539 197618 341775 197854
rect 349381 197938 349617 198174
rect 349381 197618 349617 197854
rect 357223 197938 357459 198174
rect 357223 197618 357459 197854
rect 365065 197938 365301 198174
rect 365065 197618 365301 197854
rect 375671 197938 375907 198174
rect 375671 197618 375907 197854
rect 383513 197938 383749 198174
rect 383513 197618 383749 197854
rect 391355 197938 391591 198174
rect 391355 197618 391591 197854
rect 399197 197938 399433 198174
rect 399197 197618 399433 197854
rect 409803 197938 410039 198174
rect 409803 197618 410039 197854
rect 417645 197938 417881 198174
rect 417645 197618 417881 197854
rect 425487 197938 425723 198174
rect 425487 197618 425723 197854
rect 433329 197938 433565 198174
rect 433329 197618 433565 197854
rect 443935 197938 444171 198174
rect 443935 197618 444171 197854
rect 451777 197938 452013 198174
rect 451777 197618 452013 197854
rect 459619 197938 459855 198174
rect 459619 197618 459855 197854
rect 467461 197938 467697 198174
rect 467461 197618 467697 197854
rect 478067 197938 478303 198174
rect 478067 197618 478303 197854
rect 485909 197938 486145 198174
rect 485909 197618 486145 197854
rect 493751 197938 493987 198174
rect 493751 197618 493987 197854
rect 501593 197938 501829 198174
rect 501593 197618 501829 197854
rect 512199 197938 512435 198174
rect 512199 197618 512435 197854
rect 520041 197938 520277 198174
rect 520041 197618 520277 197854
rect 527883 197938 528119 198174
rect 527883 197618 528119 197854
rect 535725 197938 535961 198174
rect 535725 197618 535961 197854
rect 546331 197938 546567 198174
rect 546331 197618 546567 197854
rect 554173 197938 554409 198174
rect 554173 197618 554409 197854
rect 562015 197938 562251 198174
rect 562015 197618 562251 197854
rect 569857 197938 570093 198174
rect 569857 197618 570093 197854
rect 337618 194218 337854 194454
rect 337618 193898 337854 194134
rect 345460 194218 345696 194454
rect 345460 193898 345696 194134
rect 353302 194218 353538 194454
rect 353302 193898 353538 194134
rect 361144 194218 361380 194454
rect 361144 193898 361380 194134
rect 371750 194218 371986 194454
rect 371750 193898 371986 194134
rect 379592 194218 379828 194454
rect 379592 193898 379828 194134
rect 387434 194218 387670 194454
rect 387434 193898 387670 194134
rect 395276 194218 395512 194454
rect 395276 193898 395512 194134
rect 405882 194218 406118 194454
rect 405882 193898 406118 194134
rect 413724 194218 413960 194454
rect 413724 193898 413960 194134
rect 421566 194218 421802 194454
rect 421566 193898 421802 194134
rect 429408 194218 429644 194454
rect 429408 193898 429644 194134
rect 440014 194218 440250 194454
rect 440014 193898 440250 194134
rect 447856 194218 448092 194454
rect 447856 193898 448092 194134
rect 455698 194218 455934 194454
rect 455698 193898 455934 194134
rect 463540 194218 463776 194454
rect 463540 193898 463776 194134
rect 474146 194218 474382 194454
rect 474146 193898 474382 194134
rect 481988 194218 482224 194454
rect 481988 193898 482224 194134
rect 489830 194218 490066 194454
rect 489830 193898 490066 194134
rect 497672 194218 497908 194454
rect 497672 193898 497908 194134
rect 508278 194218 508514 194454
rect 508278 193898 508514 194134
rect 516120 194218 516356 194454
rect 516120 193898 516356 194134
rect 523962 194218 524198 194454
rect 523962 193898 524198 194134
rect 531804 194218 532040 194454
rect 531804 193898 532040 194134
rect 542410 194218 542646 194454
rect 542410 193898 542646 194134
rect 550252 194218 550488 194454
rect 550252 193898 550488 194134
rect 558094 194218 558330 194454
rect 558094 193898 558330 194134
rect 565936 194218 566172 194454
rect 565936 193898 566172 194134
rect 337189 187938 337425 188174
rect 337189 187618 337425 187854
rect 404786 187938 405022 188174
rect 404786 187618 405022 187854
rect 472383 187938 472619 188174
rect 472383 187618 472619 187854
rect 539980 187938 540216 188174
rect 539980 187618 540216 187854
rect 303391 184218 303627 184454
rect 303391 183898 303627 184134
rect 370988 184218 371224 184454
rect 370988 183898 371224 184134
rect 438585 184218 438821 184454
rect 438585 183898 438821 184134
rect 506182 184218 506418 184454
rect 506182 183898 506418 184134
rect 307407 177643 307643 177879
rect 315249 177643 315485 177879
rect 323091 177643 323327 177879
rect 330933 177643 331169 177879
rect 303486 174218 303722 174454
rect 303486 173898 303722 174134
rect 311328 174218 311564 174454
rect 311328 173898 311564 174134
rect 319170 174218 319406 174454
rect 319170 173898 319406 174134
rect 327012 174218 327248 174454
rect 327012 173898 327248 174134
rect 307407 167938 307643 168174
rect 307407 167618 307643 167854
rect 315249 167938 315485 168174
rect 315249 167618 315485 167854
rect 323091 167938 323327 168174
rect 323091 167618 323327 167854
rect 330933 167938 331169 168174
rect 330933 167618 331169 167854
rect 303486 164218 303722 164454
rect 303486 163898 303722 164134
rect 311328 164218 311564 164454
rect 311328 163898 311564 164134
rect 319170 164218 319406 164454
rect 319170 163898 319406 164134
rect 327012 164218 327248 164454
rect 327012 163898 327248 164134
rect 293034 63935 293270 64171
rect 277674 57938 277910 58174
rect 277674 57618 277910 57854
rect 308394 57938 308630 58174
rect 308394 57618 308630 57854
rect 293034 54218 293270 54454
rect 293034 53898 293270 54134
rect 277674 47938 277910 48174
rect 277674 47618 277910 47854
rect 308394 47938 308630 48174
rect 308394 47618 308630 47854
rect 293034 44218 293270 44454
rect 293034 43898 293270 44134
rect 277674 37938 277910 38174
rect 277674 37618 277910 37854
rect 308394 37938 308630 38174
rect 308394 37618 308630 37854
rect 293034 34218 293270 34454
rect 293034 33898 293270 34134
rect 341539 177643 341775 177879
rect 349381 177643 349617 177879
rect 357223 177643 357459 177879
rect 365065 177643 365301 177879
rect 375671 177643 375907 177879
rect 383513 177643 383749 177879
rect 391355 177643 391591 177879
rect 399197 177643 399433 177879
rect 337618 174218 337854 174454
rect 337618 173898 337854 174134
rect 345460 174218 345696 174454
rect 345460 173898 345696 174134
rect 353302 174218 353538 174454
rect 353302 173898 353538 174134
rect 361144 174218 361380 174454
rect 361144 173898 361380 174134
rect 371750 174218 371986 174454
rect 371750 173898 371986 174134
rect 379592 174218 379828 174454
rect 379592 173898 379828 174134
rect 387434 174218 387670 174454
rect 387434 173898 387670 174134
rect 395276 174218 395512 174454
rect 395276 173898 395512 174134
rect 341539 167938 341775 168174
rect 341539 167618 341775 167854
rect 349381 167938 349617 168174
rect 349381 167618 349617 167854
rect 357223 167938 357459 168174
rect 357223 167618 357459 167854
rect 365065 167938 365301 168174
rect 365065 167618 365301 167854
rect 375671 167938 375907 168174
rect 375671 167618 375907 167854
rect 383513 167938 383749 168174
rect 383513 167618 383749 167854
rect 391355 167938 391591 168174
rect 391355 167618 391591 167854
rect 399197 167938 399433 168174
rect 399197 167618 399433 167854
rect 337618 164218 337854 164454
rect 337618 163898 337854 164134
rect 345460 164218 345696 164454
rect 345460 163898 345696 164134
rect 353302 164218 353538 164454
rect 353302 163898 353538 164134
rect 361144 164218 361380 164454
rect 361144 163898 361380 164134
rect 371750 164218 371986 164454
rect 371750 163898 371986 164134
rect 379592 164218 379828 164454
rect 379592 163898 379828 164134
rect 387434 164218 387670 164454
rect 387434 163898 387670 164134
rect 395276 164218 395512 164454
rect 395276 163898 395512 164134
rect 341539 157938 341775 158174
rect 341539 157618 341775 157854
rect 349381 157938 349617 158174
rect 349381 157618 349617 157854
rect 357223 157938 357459 158174
rect 357223 157618 357459 157854
rect 365065 157938 365301 158174
rect 365065 157618 365301 157854
rect 337618 154218 337854 154454
rect 337618 153898 337854 154134
rect 345460 154218 345696 154454
rect 345460 153898 345696 154134
rect 353302 154218 353538 154454
rect 353302 153898 353538 154134
rect 361144 154218 361380 154454
rect 361144 153898 361380 154134
rect 341539 147938 341775 148174
rect 341539 147618 341775 147854
rect 349381 147938 349617 148174
rect 349381 147618 349617 147854
rect 357223 147938 357459 148174
rect 357223 147618 357459 147854
rect 365065 147938 365301 148174
rect 365065 147618 365301 147854
rect 337618 144218 337854 144454
rect 337618 143898 337854 144134
rect 345460 144218 345696 144454
rect 345460 143898 345696 144134
rect 353302 144218 353538 144454
rect 353302 143898 353538 144134
rect 361144 144218 361380 144454
rect 361144 143898 361380 144134
rect 341539 137938 341775 138174
rect 341539 137618 341775 137854
rect 349381 137938 349617 138174
rect 349381 137618 349617 137854
rect 357223 137938 357459 138174
rect 357223 137618 357459 137854
rect 365065 137938 365301 138174
rect 365065 137618 365301 137854
rect 443935 177643 444171 177879
rect 451777 177643 452013 177879
rect 459619 177643 459855 177879
rect 467461 177643 467697 177879
rect 478067 177643 478303 177879
rect 485909 177643 486145 177879
rect 493751 177643 493987 177879
rect 501593 177643 501829 177879
rect 512199 177643 512435 177879
rect 520041 177643 520277 177879
rect 527883 177643 528119 177879
rect 535725 177643 535961 177879
rect 440014 174218 440250 174454
rect 440014 173898 440250 174134
rect 447856 174218 448092 174454
rect 447856 173898 448092 174134
rect 455698 174218 455934 174454
rect 455698 173898 455934 174134
rect 463540 174218 463776 174454
rect 463540 173898 463776 174134
rect 474146 174218 474382 174454
rect 474146 173898 474382 174134
rect 481988 174218 482224 174454
rect 481988 173898 482224 174134
rect 489830 174218 490066 174454
rect 489830 173898 490066 174134
rect 497672 174218 497908 174454
rect 497672 173898 497908 174134
rect 508278 174218 508514 174454
rect 508278 173898 508514 174134
rect 516120 174218 516356 174454
rect 516120 173898 516356 174134
rect 523962 174218 524198 174454
rect 523962 173898 524198 174134
rect 531804 174218 532040 174454
rect 531804 173898 532040 174134
rect 443935 167938 444171 168174
rect 443935 167618 444171 167854
rect 451777 167938 452013 168174
rect 451777 167618 452013 167854
rect 459619 167938 459855 168174
rect 459619 167618 459855 167854
rect 467461 167938 467697 168174
rect 467461 167618 467697 167854
rect 478067 167938 478303 168174
rect 478067 167618 478303 167854
rect 485909 167938 486145 168174
rect 485909 167618 486145 167854
rect 493751 167938 493987 168174
rect 493751 167618 493987 167854
rect 501593 167938 501829 168174
rect 501593 167618 501829 167854
rect 512199 167938 512435 168174
rect 512199 167618 512435 167854
rect 520041 167938 520277 168174
rect 520041 167618 520277 167854
rect 527883 167938 528119 168174
rect 527883 167618 528119 167854
rect 535725 167938 535961 168174
rect 535725 167618 535961 167854
rect 440014 164218 440250 164454
rect 440014 163898 440250 164134
rect 447856 164218 448092 164454
rect 447856 163898 448092 164134
rect 455698 164218 455934 164454
rect 455698 163898 455934 164134
rect 463540 164218 463776 164454
rect 463540 163898 463776 164134
rect 474146 164218 474382 164454
rect 474146 163898 474382 164134
rect 481988 164218 482224 164454
rect 481988 163898 482224 164134
rect 489830 164218 490066 164454
rect 489830 163898 490066 164134
rect 497672 164218 497908 164454
rect 497672 163898 497908 164134
rect 508278 164218 508514 164454
rect 508278 163898 508514 164134
rect 516120 164218 516356 164454
rect 516120 163898 516356 164134
rect 523962 164218 524198 164454
rect 523962 163898 524198 164134
rect 531804 164218 532040 164454
rect 531804 163898 532040 164134
rect 478067 157938 478303 158174
rect 478067 157618 478303 157854
rect 485909 157938 486145 158174
rect 485909 157618 486145 157854
rect 493751 157938 493987 158174
rect 493751 157618 493987 157854
rect 501593 157938 501829 158174
rect 501593 157618 501829 157854
rect 474146 154218 474382 154454
rect 474146 153898 474382 154134
rect 481988 154218 482224 154454
rect 481988 153898 482224 154134
rect 489830 154218 490066 154454
rect 489830 153898 490066 154134
rect 497672 154218 497908 154454
rect 497672 153898 497908 154134
rect 478067 147938 478303 148174
rect 478067 147618 478303 147854
rect 485909 147938 486145 148174
rect 485909 147618 486145 147854
rect 493751 147938 493987 148174
rect 493751 147618 493987 147854
rect 501593 147938 501829 148174
rect 501593 147618 501829 147854
rect 474146 144218 474382 144454
rect 474146 143898 474382 144134
rect 481988 144218 482224 144454
rect 481988 143898 482224 144134
rect 489830 144218 490066 144454
rect 489830 143898 490066 144134
rect 497672 144218 497908 144454
rect 497672 143898 497908 144134
rect 478067 137938 478303 138174
rect 478067 137618 478303 137854
rect 485909 137938 486145 138174
rect 485909 137618 486145 137854
rect 493751 137938 493987 138174
rect 493751 137618 493987 137854
rect 501593 137938 501829 138174
rect 501593 137618 501829 137854
rect 373098 127938 373334 128174
rect 373098 127618 373334 127854
rect 403818 127938 404054 128174
rect 403818 127618 404054 127854
rect 434538 127938 434774 128174
rect 434538 127618 434774 127854
rect 448186 127938 448422 128174
rect 448186 127618 448422 127854
rect 478906 127938 479142 128174
rect 478906 127618 479142 127854
rect 509626 127938 509862 128174
rect 509626 127618 509862 127854
rect 540346 127938 540582 128174
rect 540346 127618 540582 127854
rect 571066 127938 571302 128174
rect 571066 127618 571302 127854
rect 388458 124218 388694 124454
rect 388458 123898 388694 124134
rect 419178 124218 419414 124454
rect 419178 123898 419414 124134
rect 463546 124218 463782 124454
rect 463546 123898 463782 124134
rect 494266 124218 494502 124454
rect 494266 123898 494502 124134
rect 524986 124218 525222 124454
rect 524986 123898 525222 124134
rect 555706 124218 555942 124454
rect 555706 123898 555942 124134
rect 373098 117938 373334 118174
rect 373098 117618 373334 117854
rect 403818 117938 404054 118174
rect 403818 117618 404054 117854
rect 434538 117938 434774 118174
rect 434538 117618 434774 117854
rect 448186 117938 448422 118174
rect 448186 117618 448422 117854
rect 478906 117938 479142 118174
rect 478906 117618 479142 117854
rect 509626 117938 509862 118174
rect 509626 117618 509862 117854
rect 540346 117938 540582 118174
rect 540346 117618 540582 117854
rect 571066 117938 571302 118174
rect 571066 117618 571302 117854
rect 388458 114218 388694 114454
rect 388458 113898 388694 114134
rect 419178 114218 419414 114454
rect 419178 113898 419414 114134
rect 463546 114218 463782 114454
rect 463546 113898 463782 114134
rect 494266 114218 494502 114454
rect 494266 113898 494502 114134
rect 524986 114218 525222 114454
rect 524986 113898 525222 114134
rect 555706 114218 555942 114454
rect 555706 113898 555942 114134
rect 373098 107938 373334 108174
rect 373098 107618 373334 107854
rect 403818 107938 404054 108174
rect 403818 107618 404054 107854
rect 434538 107938 434774 108174
rect 434538 107618 434774 107854
rect 448186 107938 448422 108174
rect 448186 107618 448422 107854
rect 478906 107938 479142 108174
rect 478906 107618 479142 107854
rect 509626 107938 509862 108174
rect 509626 107618 509862 107854
rect 540346 107938 540582 108174
rect 540346 107618 540582 107854
rect 571066 107938 571302 108174
rect 571066 107618 571302 107854
rect 388458 104218 388694 104454
rect 388458 103898 388694 104134
rect 419178 104218 419414 104454
rect 419178 103898 419414 104134
rect 463546 104218 463782 104454
rect 463546 103898 463782 104134
rect 494266 104218 494502 104454
rect 494266 103898 494502 104134
rect 524986 104218 525222 104454
rect 524986 103898 525222 104134
rect 555706 104218 555942 104454
rect 555706 103898 555942 104134
rect 373098 97938 373334 98174
rect 373098 97618 373334 97854
rect 403818 97938 404054 98174
rect 403818 97618 404054 97854
rect 434538 97938 434774 98174
rect 434538 97618 434774 97854
rect 448186 97938 448422 98174
rect 448186 97618 448422 97854
rect 478906 97938 479142 98174
rect 478906 97618 479142 97854
rect 509626 97938 509862 98174
rect 509626 97618 509862 97854
rect 540346 97938 540582 98174
rect 540346 97618 540582 97854
rect 571066 97938 571302 98174
rect 571066 97618 571302 97854
rect 388458 94218 388694 94454
rect 388458 93898 388694 94134
rect 419178 94218 419414 94454
rect 419178 93898 419414 94134
rect 463546 94218 463782 94454
rect 463546 93898 463782 94134
rect 494266 94218 494502 94454
rect 494266 93898 494502 94134
rect 524986 94218 525222 94454
rect 524986 93898 525222 94134
rect 555706 94218 555942 94454
rect 555706 93898 555942 94134
rect 585342 667938 585578 668174
rect 585662 667938 585898 668174
rect 585342 667618 585578 667854
rect 585662 667618 585898 667854
rect 585342 657938 585578 658174
rect 585662 657938 585898 658174
rect 585342 657618 585578 657854
rect 585662 657618 585898 657854
rect 585342 647938 585578 648174
rect 585662 647938 585898 648174
rect 585342 647618 585578 647854
rect 585662 647618 585898 647854
rect 585342 637938 585578 638174
rect 585662 637938 585898 638174
rect 585342 637618 585578 637854
rect 585662 637618 585898 637854
rect 585342 627938 585578 628174
rect 585662 627938 585898 628174
rect 585342 627618 585578 627854
rect 585662 627618 585898 627854
rect 585342 617938 585578 618174
rect 585662 617938 585898 618174
rect 585342 617618 585578 617854
rect 585662 617618 585898 617854
rect 585342 607938 585578 608174
rect 585662 607938 585898 608174
rect 585342 607618 585578 607854
rect 585662 607618 585898 607854
rect 585342 597938 585578 598174
rect 585662 597938 585898 598174
rect 585342 597618 585578 597854
rect 585662 597618 585898 597854
rect 585342 587938 585578 588174
rect 585662 587938 585898 588174
rect 585342 587618 585578 587854
rect 585662 587618 585898 587854
rect 585342 577938 585578 578174
rect 585662 577938 585898 578174
rect 585342 577618 585578 577854
rect 585662 577618 585898 577854
rect 585342 567938 585578 568174
rect 585662 567938 585898 568174
rect 585342 567618 585578 567854
rect 585662 567618 585898 567854
rect 585342 557938 585578 558174
rect 585662 557938 585898 558174
rect 585342 557618 585578 557854
rect 585662 557618 585898 557854
rect 585342 547938 585578 548174
rect 585662 547938 585898 548174
rect 585342 547618 585578 547854
rect 585662 547618 585898 547854
rect 585342 537938 585578 538174
rect 585662 537938 585898 538174
rect 585342 537618 585578 537854
rect 585662 537618 585898 537854
rect 585342 527938 585578 528174
rect 585662 527938 585898 528174
rect 585342 527618 585578 527854
rect 585662 527618 585898 527854
rect 585342 517938 585578 518174
rect 585662 517938 585898 518174
rect 585342 517618 585578 517854
rect 585662 517618 585898 517854
rect 585342 507938 585578 508174
rect 585662 507938 585898 508174
rect 585342 507618 585578 507854
rect 585662 507618 585898 507854
rect 585342 497938 585578 498174
rect 585662 497938 585898 498174
rect 585342 497618 585578 497854
rect 585662 497618 585898 497854
rect 585342 487938 585578 488174
rect 585662 487938 585898 488174
rect 585342 487618 585578 487854
rect 585662 487618 585898 487854
rect 585342 477938 585578 478174
rect 585662 477938 585898 478174
rect 585342 477618 585578 477854
rect 585662 477618 585898 477854
rect 585342 467938 585578 468174
rect 585662 467938 585898 468174
rect 585342 467618 585578 467854
rect 585662 467618 585898 467854
rect 585342 457938 585578 458174
rect 585662 457938 585898 458174
rect 585342 457618 585578 457854
rect 585662 457618 585898 457854
rect 585342 447938 585578 448174
rect 585662 447938 585898 448174
rect 585342 447618 585578 447854
rect 585662 447618 585898 447854
rect 585342 437938 585578 438174
rect 585662 437938 585898 438174
rect 585342 437618 585578 437854
rect 585662 437618 585898 437854
rect 585342 427938 585578 428174
rect 585662 427938 585898 428174
rect 585342 427618 585578 427854
rect 585662 427618 585898 427854
rect 585342 417938 585578 418174
rect 585662 417938 585898 418174
rect 585342 417618 585578 417854
rect 585662 417618 585898 417854
rect 585342 407938 585578 408174
rect 585662 407938 585898 408174
rect 585342 407618 585578 407854
rect 585662 407618 585898 407854
rect 585342 397938 585578 398174
rect 585662 397938 585898 398174
rect 585342 397618 585578 397854
rect 585662 397618 585898 397854
rect 585342 387938 585578 388174
rect 585662 387938 585898 388174
rect 585342 387618 585578 387854
rect 585662 387618 585898 387854
rect 585342 377938 585578 378174
rect 585662 377938 585898 378174
rect 585342 377618 585578 377854
rect 585662 377618 585898 377854
rect 585342 367938 585578 368174
rect 585662 367938 585898 368174
rect 585342 367618 585578 367854
rect 585662 367618 585898 367854
rect 585342 357938 585578 358174
rect 585662 357938 585898 358174
rect 585342 357618 585578 357854
rect 585662 357618 585898 357854
rect 585342 347938 585578 348174
rect 585662 347938 585898 348174
rect 585342 347618 585578 347854
rect 585662 347618 585898 347854
rect 585342 337938 585578 338174
rect 585662 337938 585898 338174
rect 585342 337618 585578 337854
rect 585662 337618 585898 337854
rect 585342 327938 585578 328174
rect 585662 327938 585898 328174
rect 585342 327618 585578 327854
rect 585662 327618 585898 327854
rect 585342 317938 585578 318174
rect 585662 317938 585898 318174
rect 585342 317618 585578 317854
rect 585662 317618 585898 317854
rect 585342 307938 585578 308174
rect 585662 307938 585898 308174
rect 585342 307618 585578 307854
rect 585662 307618 585898 307854
rect 585342 297938 585578 298174
rect 585662 297938 585898 298174
rect 585342 297618 585578 297854
rect 585662 297618 585898 297854
rect 585342 287938 585578 288174
rect 585662 287938 585898 288174
rect 585342 287618 585578 287854
rect 585662 287618 585898 287854
rect 585342 277938 585578 278174
rect 585662 277938 585898 278174
rect 585342 277618 585578 277854
rect 585662 277618 585898 277854
rect 585342 267938 585578 268174
rect 585662 267938 585898 268174
rect 585342 267618 585578 267854
rect 585662 267618 585898 267854
rect 585342 257938 585578 258174
rect 585662 257938 585898 258174
rect 585342 257618 585578 257854
rect 585662 257618 585898 257854
rect 585342 247938 585578 248174
rect 585662 247938 585898 248174
rect 585342 247618 585578 247854
rect 585662 247618 585898 247854
rect 585342 237938 585578 238174
rect 585662 237938 585898 238174
rect 585342 237618 585578 237854
rect 585662 237618 585898 237854
rect 585342 227938 585578 228174
rect 585662 227938 585898 228174
rect 585342 227618 585578 227854
rect 585662 227618 585898 227854
rect 585342 217938 585578 218174
rect 585662 217938 585898 218174
rect 585342 217618 585578 217854
rect 585662 217618 585898 217854
rect 585342 207938 585578 208174
rect 585662 207938 585898 208174
rect 585342 207618 585578 207854
rect 585662 207618 585898 207854
rect 585342 197938 585578 198174
rect 585662 197938 585898 198174
rect 585342 197618 585578 197854
rect 585662 197618 585898 197854
rect 585342 187938 585578 188174
rect 585662 187938 585898 188174
rect 585342 187618 585578 187854
rect 585662 187618 585898 187854
rect 585342 177938 585578 178174
rect 585662 177938 585898 178174
rect 585342 177618 585578 177854
rect 585662 177618 585898 177854
rect 585342 167938 585578 168174
rect 585662 167938 585898 168174
rect 585342 167618 585578 167854
rect 585662 167618 585898 167854
rect 585342 157938 585578 158174
rect 585662 157938 585898 158174
rect 585342 157618 585578 157854
rect 585662 157618 585898 157854
rect 585342 147938 585578 148174
rect 585662 147938 585898 148174
rect 585342 147618 585578 147854
rect 585662 147618 585898 147854
rect 585342 137938 585578 138174
rect 585662 137938 585898 138174
rect 585342 137618 585578 137854
rect 585662 137618 585898 137854
rect 585342 127938 585578 128174
rect 585662 127938 585898 128174
rect 585342 127618 585578 127854
rect 585662 127618 585898 127854
rect 585342 117938 585578 118174
rect 585662 117938 585898 118174
rect 585342 117618 585578 117854
rect 585662 117618 585898 117854
rect 585342 107938 585578 108174
rect 585662 107938 585898 108174
rect 585342 107618 585578 107854
rect 585662 107618 585898 107854
rect 585342 97938 585578 98174
rect 585662 97938 585898 98174
rect 585342 97618 585578 97854
rect 585662 97618 585898 97854
rect 585342 87938 585578 88174
rect 585662 87938 585898 88174
rect 585342 87618 585578 87854
rect 585662 87618 585898 87854
rect 585342 77938 585578 78174
rect 585662 77938 585898 78174
rect 585342 77618 585578 77854
rect 585662 77618 585898 77854
rect 585342 67938 585578 68174
rect 585662 67938 585898 68174
rect 585342 67618 585578 67854
rect 585662 67618 585898 67854
rect 585342 57938 585578 58174
rect 585662 57938 585898 58174
rect 585342 57618 585578 57854
rect 585662 57618 585898 57854
rect 585342 47938 585578 48174
rect 585662 47938 585898 48174
rect 585342 47618 585578 47854
rect 585662 47618 585898 47854
rect 585342 37938 585578 38174
rect 585662 37938 585898 38174
rect 585342 37618 585578 37854
rect 585662 37618 585898 37854
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 694218 586538 694454
rect 586622 694218 586858 694454
rect 586302 693898 586538 694134
rect 586622 693898 586858 694134
rect 586302 684218 586538 684454
rect 586622 684218 586858 684454
rect 586302 683898 586538 684134
rect 586622 683898 586858 684134
rect 586302 674218 586538 674454
rect 586622 674218 586858 674454
rect 586302 673898 586538 674134
rect 586622 673898 586858 674134
rect 586302 664218 586538 664454
rect 586622 664218 586858 664454
rect 586302 663898 586538 664134
rect 586622 663898 586858 664134
rect 586302 654218 586538 654454
rect 586622 654218 586858 654454
rect 586302 653898 586538 654134
rect 586622 653898 586858 654134
rect 586302 644218 586538 644454
rect 586622 644218 586858 644454
rect 586302 643898 586538 644134
rect 586622 643898 586858 644134
rect 586302 634218 586538 634454
rect 586622 634218 586858 634454
rect 586302 633898 586538 634134
rect 586622 633898 586858 634134
rect 586302 624218 586538 624454
rect 586622 624218 586858 624454
rect 586302 623898 586538 624134
rect 586622 623898 586858 624134
rect 586302 614218 586538 614454
rect 586622 614218 586858 614454
rect 586302 613898 586538 614134
rect 586622 613898 586858 614134
rect 586302 604218 586538 604454
rect 586622 604218 586858 604454
rect 586302 603898 586538 604134
rect 586622 603898 586858 604134
rect 586302 594218 586538 594454
rect 586622 594218 586858 594454
rect 586302 593898 586538 594134
rect 586622 593898 586858 594134
rect 586302 584218 586538 584454
rect 586622 584218 586858 584454
rect 586302 583898 586538 584134
rect 586622 583898 586858 584134
rect 586302 574218 586538 574454
rect 586622 574218 586858 574454
rect 586302 573898 586538 574134
rect 586622 573898 586858 574134
rect 586302 564218 586538 564454
rect 586622 564218 586858 564454
rect 586302 563898 586538 564134
rect 586622 563898 586858 564134
rect 586302 554218 586538 554454
rect 586622 554218 586858 554454
rect 586302 553898 586538 554134
rect 586622 553898 586858 554134
rect 586302 544218 586538 544454
rect 586622 544218 586858 544454
rect 586302 543898 586538 544134
rect 586622 543898 586858 544134
rect 586302 534218 586538 534454
rect 586622 534218 586858 534454
rect 586302 533898 586538 534134
rect 586622 533898 586858 534134
rect 586302 524218 586538 524454
rect 586622 524218 586858 524454
rect 586302 523898 586538 524134
rect 586622 523898 586858 524134
rect 586302 514218 586538 514454
rect 586622 514218 586858 514454
rect 586302 513898 586538 514134
rect 586622 513898 586858 514134
rect 586302 504218 586538 504454
rect 586622 504218 586858 504454
rect 586302 503898 586538 504134
rect 586622 503898 586858 504134
rect 586302 494218 586538 494454
rect 586622 494218 586858 494454
rect 586302 493898 586538 494134
rect 586622 493898 586858 494134
rect 586302 484218 586538 484454
rect 586622 484218 586858 484454
rect 586302 483898 586538 484134
rect 586622 483898 586858 484134
rect 586302 474218 586538 474454
rect 586622 474218 586858 474454
rect 586302 473898 586538 474134
rect 586622 473898 586858 474134
rect 586302 464218 586538 464454
rect 586622 464218 586858 464454
rect 586302 463898 586538 464134
rect 586622 463898 586858 464134
rect 586302 454218 586538 454454
rect 586622 454218 586858 454454
rect 586302 453898 586538 454134
rect 586622 453898 586858 454134
rect 586302 444218 586538 444454
rect 586622 444218 586858 444454
rect 586302 443898 586538 444134
rect 586622 443898 586858 444134
rect 586302 434218 586538 434454
rect 586622 434218 586858 434454
rect 586302 433898 586538 434134
rect 586622 433898 586858 434134
rect 586302 424218 586538 424454
rect 586622 424218 586858 424454
rect 586302 423898 586538 424134
rect 586622 423898 586858 424134
rect 586302 414218 586538 414454
rect 586622 414218 586858 414454
rect 586302 413898 586538 414134
rect 586622 413898 586858 414134
rect 586302 404218 586538 404454
rect 586622 404218 586858 404454
rect 586302 403898 586538 404134
rect 586622 403898 586858 404134
rect 586302 394218 586538 394454
rect 586622 394218 586858 394454
rect 586302 393898 586538 394134
rect 586622 393898 586858 394134
rect 586302 384218 586538 384454
rect 586622 384218 586858 384454
rect 586302 383898 586538 384134
rect 586622 383898 586858 384134
rect 586302 374218 586538 374454
rect 586622 374218 586858 374454
rect 586302 373898 586538 374134
rect 586622 373898 586858 374134
rect 586302 364218 586538 364454
rect 586622 364218 586858 364454
rect 586302 363898 586538 364134
rect 586622 363898 586858 364134
rect 586302 354218 586538 354454
rect 586622 354218 586858 354454
rect 586302 353898 586538 354134
rect 586622 353898 586858 354134
rect 586302 344218 586538 344454
rect 586622 344218 586858 344454
rect 586302 343898 586538 344134
rect 586622 343898 586858 344134
rect 586302 334218 586538 334454
rect 586622 334218 586858 334454
rect 586302 333898 586538 334134
rect 586622 333898 586858 334134
rect 586302 324218 586538 324454
rect 586622 324218 586858 324454
rect 586302 323898 586538 324134
rect 586622 323898 586858 324134
rect 586302 314218 586538 314454
rect 586622 314218 586858 314454
rect 586302 313898 586538 314134
rect 586622 313898 586858 314134
rect 586302 304218 586538 304454
rect 586622 304218 586858 304454
rect 586302 303898 586538 304134
rect 586622 303898 586858 304134
rect 586302 294218 586538 294454
rect 586622 294218 586858 294454
rect 586302 293898 586538 294134
rect 586622 293898 586858 294134
rect 586302 284218 586538 284454
rect 586622 284218 586858 284454
rect 586302 283898 586538 284134
rect 586622 283898 586858 284134
rect 586302 274218 586538 274454
rect 586622 274218 586858 274454
rect 586302 273898 586538 274134
rect 586622 273898 586858 274134
rect 586302 264218 586538 264454
rect 586622 264218 586858 264454
rect 586302 263898 586538 264134
rect 586622 263898 586858 264134
rect 586302 254218 586538 254454
rect 586622 254218 586858 254454
rect 586302 253898 586538 254134
rect 586622 253898 586858 254134
rect 586302 244218 586538 244454
rect 586622 244218 586858 244454
rect 586302 243898 586538 244134
rect 586622 243898 586858 244134
rect 586302 234218 586538 234454
rect 586622 234218 586858 234454
rect 586302 233898 586538 234134
rect 586622 233898 586858 234134
rect 586302 224218 586538 224454
rect 586622 224218 586858 224454
rect 586302 223898 586538 224134
rect 586622 223898 586858 224134
rect 586302 214218 586538 214454
rect 586622 214218 586858 214454
rect 586302 213898 586538 214134
rect 586622 213898 586858 214134
rect 586302 204218 586538 204454
rect 586622 204218 586858 204454
rect 586302 203898 586538 204134
rect 586622 203898 586858 204134
rect 586302 194218 586538 194454
rect 586622 194218 586858 194454
rect 586302 193898 586538 194134
rect 586622 193898 586858 194134
rect 586302 184218 586538 184454
rect 586622 184218 586858 184454
rect 586302 183898 586538 184134
rect 586622 183898 586858 184134
rect 586302 174218 586538 174454
rect 586622 174218 586858 174454
rect 586302 173898 586538 174134
rect 586622 173898 586858 174134
rect 586302 164218 586538 164454
rect 586622 164218 586858 164454
rect 586302 163898 586538 164134
rect 586622 163898 586858 164134
rect 586302 154218 586538 154454
rect 586622 154218 586858 154454
rect 586302 153898 586538 154134
rect 586622 153898 586858 154134
rect 586302 144218 586538 144454
rect 586622 144218 586858 144454
rect 586302 143898 586538 144134
rect 586622 143898 586858 144134
rect 586302 134218 586538 134454
rect 586622 134218 586858 134454
rect 586302 133898 586538 134134
rect 586622 133898 586858 134134
rect 586302 124218 586538 124454
rect 586622 124218 586858 124454
rect 586302 123898 586538 124134
rect 586622 123898 586858 124134
rect 586302 114218 586538 114454
rect 586622 114218 586858 114454
rect 586302 113898 586538 114134
rect 586622 113898 586858 114134
rect 586302 104218 586538 104454
rect 586622 104218 586858 104454
rect 586302 103898 586538 104134
rect 586622 103898 586858 104134
rect 586302 94218 586538 94454
rect 586622 94218 586858 94454
rect 586302 93898 586538 94134
rect 586622 93898 586858 94134
rect 586302 84218 586538 84454
rect 586622 84218 586858 84454
rect 586302 83898 586538 84134
rect 586622 83898 586858 84134
rect 586302 74218 586538 74454
rect 586622 74218 586858 74454
rect 586302 73898 586538 74134
rect 586622 73898 586858 74134
rect 586302 64218 586538 64454
rect 586622 64218 586858 64454
rect 586302 63898 586538 64134
rect 586622 63898 586858 64134
rect 586302 54218 586538 54454
rect 586622 54218 586858 54454
rect 586302 53898 586538 54134
rect 586622 53898 586858 54134
rect 586302 44218 586538 44454
rect 586622 44218 586858 44454
rect 586302 43898 586538 44134
rect 586622 43898 586858 44134
rect 586302 34218 586538 34454
rect 586622 34218 586858 34454
rect 586302 33898 586538 34134
rect 586622 33898 586858 34134
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698174 592650 698206
rect -8726 697938 -1974 698174
rect -1738 697938 -1654 698174
rect -1418 697938 585342 698174
rect 585578 697938 585662 698174
rect 585898 697938 592650 698174
rect -8726 697854 592650 697938
rect -8726 697618 -1974 697854
rect -1738 697618 -1654 697854
rect -1418 697618 585342 697854
rect 585578 697618 585662 697854
rect 585898 697618 592650 697854
rect -8726 697586 592650 697618
rect -8726 694454 592650 694486
rect -8726 694218 -2934 694454
rect -2698 694218 -2614 694454
rect -2378 694218 586302 694454
rect 586538 694218 586622 694454
rect 586858 694218 592650 694454
rect -8726 694134 592650 694218
rect -8726 693898 -2934 694134
rect -2698 693898 -2614 694134
rect -2378 693898 586302 694134
rect 586538 693898 586622 694134
rect 586858 693898 592650 694134
rect -8726 693866 592650 693898
rect -8726 688174 592650 688206
rect -8726 687938 -1974 688174
rect -1738 687938 -1654 688174
rect -1418 687938 585342 688174
rect 585578 687938 585662 688174
rect 585898 687938 592650 688174
rect -8726 687854 592650 687938
rect -8726 687618 -1974 687854
rect -1738 687618 -1654 687854
rect -1418 687618 585342 687854
rect 585578 687618 585662 687854
rect 585898 687618 592650 687854
rect -8726 687586 592650 687618
rect -8726 684454 592650 684486
rect -8726 684218 -2934 684454
rect -2698 684218 -2614 684454
rect -2378 684218 586302 684454
rect 586538 684218 586622 684454
rect 586858 684218 592650 684454
rect -8726 684134 592650 684218
rect -8726 683898 -2934 684134
rect -2698 683898 -2614 684134
rect -2378 683898 586302 684134
rect 586538 683898 586622 684134
rect 586858 683898 592650 684134
rect -8726 683866 592650 683898
rect -8726 678174 592650 678206
rect -8726 677938 -1974 678174
rect -1738 677938 -1654 678174
rect -1418 677938 585342 678174
rect 585578 677938 585662 678174
rect 585898 677938 592650 678174
rect -8726 677854 592650 677938
rect -8726 677618 -1974 677854
rect -1738 677618 -1654 677854
rect -1418 677618 585342 677854
rect 585578 677618 585662 677854
rect 585898 677618 592650 677854
rect -8726 677586 592650 677618
rect -8726 674454 592650 674486
rect -8726 674218 -2934 674454
rect -2698 674218 -2614 674454
rect -2378 674218 586302 674454
rect 586538 674218 586622 674454
rect 586858 674218 592650 674454
rect -8726 674134 592650 674218
rect -8726 673898 -2934 674134
rect -2698 673898 -2614 674134
rect -2378 673898 586302 674134
rect 586538 673898 586622 674134
rect 586858 673898 592650 674134
rect -8726 673866 592650 673898
rect -8726 668174 592650 668206
rect -8726 667938 -1974 668174
rect -1738 667938 -1654 668174
rect -1418 667938 585342 668174
rect 585578 667938 585662 668174
rect 585898 667938 592650 668174
rect -8726 667854 592650 667938
rect -8726 667618 -1974 667854
rect -1738 667618 -1654 667854
rect -1418 667618 585342 667854
rect 585578 667618 585662 667854
rect 585898 667618 592650 667854
rect -8726 667586 592650 667618
rect -8726 664454 592650 664486
rect -8726 664218 -2934 664454
rect -2698 664218 -2614 664454
rect -2378 664218 586302 664454
rect 586538 664218 586622 664454
rect 586858 664218 592650 664454
rect -8726 664134 592650 664218
rect -8726 663898 -2934 664134
rect -2698 663898 -2614 664134
rect -2378 663898 586302 664134
rect 586538 663898 586622 664134
rect 586858 663898 592650 664134
rect -8726 663866 592650 663898
rect -8726 658174 592650 658206
rect -8726 657938 -1974 658174
rect -1738 657938 -1654 658174
rect -1418 657938 585342 658174
rect 585578 657938 585662 658174
rect 585898 657938 592650 658174
rect -8726 657854 592650 657938
rect -8726 657618 -1974 657854
rect -1738 657618 -1654 657854
rect -1418 657618 585342 657854
rect 585578 657618 585662 657854
rect 585898 657618 592650 657854
rect -8726 657586 592650 657618
rect -8726 654454 592650 654486
rect -8726 654218 -2934 654454
rect -2698 654218 -2614 654454
rect -2378 654218 586302 654454
rect 586538 654218 586622 654454
rect 586858 654218 592650 654454
rect -8726 654134 592650 654218
rect -8726 653898 -2934 654134
rect -2698 653898 -2614 654134
rect -2378 653898 586302 654134
rect 586538 653898 586622 654134
rect 586858 653898 592650 654134
rect -8726 653866 592650 653898
rect -8726 648174 592650 648206
rect -8726 647938 -1974 648174
rect -1738 647938 -1654 648174
rect -1418 647938 585342 648174
rect 585578 647938 585662 648174
rect 585898 647938 592650 648174
rect -8726 647854 592650 647938
rect -8726 647618 -1974 647854
rect -1738 647618 -1654 647854
rect -1418 647618 585342 647854
rect 585578 647618 585662 647854
rect 585898 647618 592650 647854
rect -8726 647586 592650 647618
rect -8726 644454 592650 644486
rect -8726 644218 -2934 644454
rect -2698 644218 -2614 644454
rect -2378 644218 586302 644454
rect 586538 644218 586622 644454
rect 586858 644218 592650 644454
rect -8726 644134 592650 644218
rect -8726 643898 -2934 644134
rect -2698 643898 -2614 644134
rect -2378 643898 586302 644134
rect 586538 643898 586622 644134
rect 586858 643898 592650 644134
rect -8726 643866 592650 643898
rect -8726 638174 592650 638206
rect -8726 637938 -1974 638174
rect -1738 637938 -1654 638174
rect -1418 637938 585342 638174
rect 585578 637938 585662 638174
rect 585898 637938 592650 638174
rect -8726 637854 592650 637938
rect -8726 637618 -1974 637854
rect -1738 637618 -1654 637854
rect -1418 637618 585342 637854
rect 585578 637618 585662 637854
rect 585898 637618 592650 637854
rect -8726 637586 592650 637618
rect -8726 634454 592650 634486
rect -8726 634218 -2934 634454
rect -2698 634218 -2614 634454
rect -2378 634218 586302 634454
rect 586538 634218 586622 634454
rect 586858 634218 592650 634454
rect -8726 634134 592650 634218
rect -8726 633898 -2934 634134
rect -2698 633898 -2614 634134
rect -2378 633898 586302 634134
rect 586538 633898 586622 634134
rect 586858 633898 592650 634134
rect -8726 633866 592650 633898
rect -8726 628174 592650 628206
rect -8726 627938 -1974 628174
rect -1738 627938 -1654 628174
rect -1418 627938 585342 628174
rect 585578 627938 585662 628174
rect 585898 627938 592650 628174
rect -8726 627854 592650 627938
rect -8726 627618 -1974 627854
rect -1738 627618 -1654 627854
rect -1418 627618 585342 627854
rect 585578 627618 585662 627854
rect 585898 627618 592650 627854
rect -8726 627586 592650 627618
rect -8726 624454 592650 624486
rect -8726 624218 -2934 624454
rect -2698 624218 -2614 624454
rect -2378 624218 586302 624454
rect 586538 624218 586622 624454
rect 586858 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -2934 624134
rect -2698 623898 -2614 624134
rect -2378 623898 586302 624134
rect 586538 623898 586622 624134
rect 586858 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 618174 592650 618206
rect -8726 617938 -1974 618174
rect -1738 617938 -1654 618174
rect -1418 617938 585342 618174
rect 585578 617938 585662 618174
rect 585898 617938 592650 618174
rect -8726 617854 592650 617938
rect -8726 617618 -1974 617854
rect -1738 617618 -1654 617854
rect -1418 617618 585342 617854
rect 585578 617618 585662 617854
rect 585898 617618 592650 617854
rect -8726 617586 592650 617618
rect -8726 614454 592650 614486
rect -8726 614218 -2934 614454
rect -2698 614218 -2614 614454
rect -2378 614218 586302 614454
rect 586538 614218 586622 614454
rect 586858 614218 592650 614454
rect -8726 614134 592650 614218
rect -8726 613898 -2934 614134
rect -2698 613898 -2614 614134
rect -2378 613898 586302 614134
rect 586538 613898 586622 614134
rect 586858 613898 592650 614134
rect -8726 613866 592650 613898
rect -8726 608174 592650 608206
rect -8726 607938 -1974 608174
rect -1738 607938 -1654 608174
rect -1418 607938 585342 608174
rect 585578 607938 585662 608174
rect 585898 607938 592650 608174
rect -8726 607854 592650 607938
rect -8726 607618 -1974 607854
rect -1738 607618 -1654 607854
rect -1418 607618 585342 607854
rect 585578 607618 585662 607854
rect 585898 607618 592650 607854
rect -8726 607586 592650 607618
rect -8726 604454 592650 604486
rect -8726 604218 -2934 604454
rect -2698 604218 -2614 604454
rect -2378 604218 586302 604454
rect 586538 604218 586622 604454
rect 586858 604218 592650 604454
rect -8726 604134 592650 604218
rect -8726 603898 -2934 604134
rect -2698 603898 -2614 604134
rect -2378 603898 586302 604134
rect 586538 603898 586622 604134
rect 586858 603898 592650 604134
rect -8726 603866 592650 603898
rect -8726 598174 592650 598206
rect -8726 597938 -1974 598174
rect -1738 597938 -1654 598174
rect -1418 597938 585342 598174
rect 585578 597938 585662 598174
rect 585898 597938 592650 598174
rect -8726 597854 592650 597938
rect -8726 597618 -1974 597854
rect -1738 597618 -1654 597854
rect -1418 597618 585342 597854
rect 585578 597618 585662 597854
rect 585898 597618 592650 597854
rect -8726 597586 592650 597618
rect -8726 594454 592650 594486
rect -8726 594218 -2934 594454
rect -2698 594218 -2614 594454
rect -2378 594218 586302 594454
rect 586538 594218 586622 594454
rect 586858 594218 592650 594454
rect -8726 594134 592650 594218
rect -8726 593898 -2934 594134
rect -2698 593898 -2614 594134
rect -2378 593898 586302 594134
rect 586538 593898 586622 594134
rect 586858 593898 592650 594134
rect -8726 593866 592650 593898
rect -8726 588174 592650 588206
rect -8726 587938 -1974 588174
rect -1738 587938 -1654 588174
rect -1418 587938 585342 588174
rect 585578 587938 585662 588174
rect 585898 587938 592650 588174
rect -8726 587854 592650 587938
rect -8726 587618 -1974 587854
rect -1738 587618 -1654 587854
rect -1418 587618 585342 587854
rect 585578 587618 585662 587854
rect 585898 587618 592650 587854
rect -8726 587586 592650 587618
rect -8726 584454 592650 584486
rect -8726 584218 -2934 584454
rect -2698 584218 -2614 584454
rect -2378 584218 586302 584454
rect 586538 584218 586622 584454
rect 586858 584218 592650 584454
rect -8726 584134 592650 584218
rect -8726 583898 -2934 584134
rect -2698 583898 -2614 584134
rect -2378 583898 586302 584134
rect 586538 583898 586622 584134
rect 586858 583898 592650 584134
rect -8726 583866 592650 583898
rect -8726 578174 592650 578206
rect -8726 577938 -1974 578174
rect -1738 577938 -1654 578174
rect -1418 577938 585342 578174
rect 585578 577938 585662 578174
rect 585898 577938 592650 578174
rect -8726 577854 592650 577938
rect -8726 577618 -1974 577854
rect -1738 577618 -1654 577854
rect -1418 577618 585342 577854
rect 585578 577618 585662 577854
rect 585898 577618 592650 577854
rect -8726 577586 592650 577618
rect -8726 574454 592650 574486
rect -8726 574218 -2934 574454
rect -2698 574218 -2614 574454
rect -2378 574218 586302 574454
rect 586538 574218 586622 574454
rect 586858 574218 592650 574454
rect -8726 574134 592650 574218
rect -8726 573898 -2934 574134
rect -2698 573898 -2614 574134
rect -2378 573898 586302 574134
rect 586538 573898 586622 574134
rect 586858 573898 592650 574134
rect -8726 573866 592650 573898
rect -8726 568174 592650 568206
rect -8726 567938 -1974 568174
rect -1738 567938 -1654 568174
rect -1418 567938 585342 568174
rect 585578 567938 585662 568174
rect 585898 567938 592650 568174
rect -8726 567854 592650 567938
rect -8726 567618 -1974 567854
rect -1738 567618 -1654 567854
rect -1418 567618 585342 567854
rect 585578 567618 585662 567854
rect 585898 567618 592650 567854
rect -8726 567586 592650 567618
rect -8726 564454 592650 564486
rect -8726 564218 -2934 564454
rect -2698 564218 -2614 564454
rect -2378 564218 586302 564454
rect 586538 564218 586622 564454
rect 586858 564218 592650 564454
rect -8726 564134 592650 564218
rect -8726 563898 -2934 564134
rect -2698 563898 -2614 564134
rect -2378 563898 586302 564134
rect 586538 563898 586622 564134
rect 586858 563898 592650 564134
rect -8726 563866 592650 563898
rect -8726 558174 592650 558206
rect -8726 557938 -1974 558174
rect -1738 557938 -1654 558174
rect -1418 557938 585342 558174
rect 585578 557938 585662 558174
rect 585898 557938 592650 558174
rect -8726 557854 592650 557938
rect -8726 557618 -1974 557854
rect -1738 557618 -1654 557854
rect -1418 557618 585342 557854
rect 585578 557618 585662 557854
rect 585898 557618 592650 557854
rect -8726 557586 592650 557618
rect -8726 554454 592650 554486
rect -8726 554218 -2934 554454
rect -2698 554218 -2614 554454
rect -2378 554218 586302 554454
rect 586538 554218 586622 554454
rect 586858 554218 592650 554454
rect -8726 554134 592650 554218
rect -8726 553898 -2934 554134
rect -2698 553898 -2614 554134
rect -2378 553898 586302 554134
rect 586538 553898 586622 554134
rect 586858 553898 592650 554134
rect -8726 553866 592650 553898
rect -8726 548174 592650 548206
rect -8726 547938 -1974 548174
rect -1738 547938 -1654 548174
rect -1418 547938 585342 548174
rect 585578 547938 585662 548174
rect 585898 547938 592650 548174
rect -8726 547854 592650 547938
rect -8726 547618 -1974 547854
rect -1738 547618 -1654 547854
rect -1418 547618 585342 547854
rect 585578 547618 585662 547854
rect 585898 547618 592650 547854
rect -8726 547586 592650 547618
rect -8726 544454 592650 544486
rect -8726 544218 -2934 544454
rect -2698 544218 -2614 544454
rect -2378 544218 586302 544454
rect 586538 544218 586622 544454
rect 586858 544218 592650 544454
rect -8726 544134 592650 544218
rect -8726 543898 -2934 544134
rect -2698 543898 -2614 544134
rect -2378 543898 586302 544134
rect 586538 543898 586622 544134
rect 586858 543898 592650 544134
rect -8726 543866 592650 543898
rect -8726 538174 592650 538206
rect -8726 537938 -1974 538174
rect -1738 537938 -1654 538174
rect -1418 537938 585342 538174
rect 585578 537938 585662 538174
rect 585898 537938 592650 538174
rect -8726 537854 592650 537938
rect -8726 537618 -1974 537854
rect -1738 537618 -1654 537854
rect -1418 537618 585342 537854
rect 585578 537618 585662 537854
rect 585898 537618 592650 537854
rect -8726 537586 592650 537618
rect -8726 534454 592650 534486
rect -8726 534218 -2934 534454
rect -2698 534218 -2614 534454
rect -2378 534218 586302 534454
rect 586538 534218 586622 534454
rect 586858 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -2934 534134
rect -2698 533898 -2614 534134
rect -2378 533898 586302 534134
rect 586538 533898 586622 534134
rect 586858 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 528174 592650 528206
rect -8726 527938 -1974 528174
rect -1738 527938 -1654 528174
rect -1418 527938 585342 528174
rect 585578 527938 585662 528174
rect 585898 527938 592650 528174
rect -8726 527854 592650 527938
rect -8726 527618 -1974 527854
rect -1738 527618 -1654 527854
rect -1418 527618 585342 527854
rect 585578 527618 585662 527854
rect 585898 527618 592650 527854
rect -8726 527586 592650 527618
rect -8726 524454 592650 524486
rect -8726 524218 -2934 524454
rect -2698 524218 -2614 524454
rect -2378 524218 586302 524454
rect 586538 524218 586622 524454
rect 586858 524218 592650 524454
rect -8726 524134 592650 524218
rect -8726 523898 -2934 524134
rect -2698 523898 -2614 524134
rect -2378 523898 586302 524134
rect 586538 523898 586622 524134
rect 586858 523898 592650 524134
rect -8726 523866 592650 523898
rect -8726 518174 592650 518206
rect -8726 517938 -1974 518174
rect -1738 517938 -1654 518174
rect -1418 517938 585342 518174
rect 585578 517938 585662 518174
rect 585898 517938 592650 518174
rect -8726 517854 592650 517938
rect -8726 517618 -1974 517854
rect -1738 517618 -1654 517854
rect -1418 517618 585342 517854
rect 585578 517618 585662 517854
rect 585898 517618 592650 517854
rect -8726 517586 592650 517618
rect -8726 514454 592650 514486
rect -8726 514218 -2934 514454
rect -2698 514218 -2614 514454
rect -2378 514218 586302 514454
rect 586538 514218 586622 514454
rect 586858 514218 592650 514454
rect -8726 514134 592650 514218
rect -8726 513898 -2934 514134
rect -2698 513898 -2614 514134
rect -2378 513898 586302 514134
rect 586538 513898 586622 514134
rect 586858 513898 592650 514134
rect -8726 513866 592650 513898
rect -8726 508174 592650 508206
rect -8726 507938 -1974 508174
rect -1738 507938 -1654 508174
rect -1418 507938 585342 508174
rect 585578 507938 585662 508174
rect 585898 507938 592650 508174
rect -8726 507854 592650 507938
rect -8726 507618 -1974 507854
rect -1738 507618 -1654 507854
rect -1418 507618 585342 507854
rect 585578 507618 585662 507854
rect 585898 507618 592650 507854
rect -8726 507586 592650 507618
rect -8726 504454 592650 504486
rect -8726 504218 -2934 504454
rect -2698 504218 -2614 504454
rect -2378 504218 586302 504454
rect 586538 504218 586622 504454
rect 586858 504218 592650 504454
rect -8726 504134 592650 504218
rect -8726 503898 -2934 504134
rect -2698 503898 -2614 504134
rect -2378 503898 586302 504134
rect 586538 503898 586622 504134
rect 586858 503898 592650 504134
rect -8726 503866 592650 503898
rect -8726 498174 592650 498206
rect -8726 497938 -1974 498174
rect -1738 497938 -1654 498174
rect -1418 497938 585342 498174
rect 585578 497938 585662 498174
rect 585898 497938 592650 498174
rect -8726 497854 592650 497938
rect -8726 497618 -1974 497854
rect -1738 497618 -1654 497854
rect -1418 497618 585342 497854
rect 585578 497618 585662 497854
rect 585898 497618 592650 497854
rect -8726 497586 592650 497618
rect -8726 494454 592650 494486
rect -8726 494218 -2934 494454
rect -2698 494218 -2614 494454
rect -2378 494218 586302 494454
rect 586538 494218 586622 494454
rect 586858 494218 592650 494454
rect -8726 494134 592650 494218
rect -8726 493898 -2934 494134
rect -2698 493898 -2614 494134
rect -2378 493898 586302 494134
rect 586538 493898 586622 494134
rect 586858 493898 592650 494134
rect -8726 493866 592650 493898
rect -8726 488174 592650 488206
rect -8726 487938 -1974 488174
rect -1738 487938 -1654 488174
rect -1418 487938 585342 488174
rect 585578 487938 585662 488174
rect 585898 487938 592650 488174
rect -8726 487854 592650 487938
rect -8726 487618 -1974 487854
rect -1738 487618 -1654 487854
rect -1418 487618 585342 487854
rect 585578 487618 585662 487854
rect 585898 487618 592650 487854
rect -8726 487586 592650 487618
rect -8726 484454 592650 484486
rect -8726 484218 -2934 484454
rect -2698 484218 -2614 484454
rect -2378 484218 586302 484454
rect 586538 484218 586622 484454
rect 586858 484218 592650 484454
rect -8726 484134 592650 484218
rect -8726 483898 -2934 484134
rect -2698 483898 -2614 484134
rect -2378 483898 586302 484134
rect 586538 483898 586622 484134
rect 586858 483898 592650 484134
rect -8726 483866 592650 483898
rect -8726 478174 592650 478206
rect -8726 477938 -1974 478174
rect -1738 477938 -1654 478174
rect -1418 477938 585342 478174
rect 585578 477938 585662 478174
rect 585898 477938 592650 478174
rect -8726 477854 592650 477938
rect -8726 477618 -1974 477854
rect -1738 477618 -1654 477854
rect -1418 477618 585342 477854
rect 585578 477618 585662 477854
rect 585898 477618 592650 477854
rect -8726 477586 592650 477618
rect -8726 474454 592650 474486
rect -8726 474218 -2934 474454
rect -2698 474218 -2614 474454
rect -2378 474218 586302 474454
rect 586538 474218 586622 474454
rect 586858 474218 592650 474454
rect -8726 474134 592650 474218
rect -8726 473898 -2934 474134
rect -2698 473898 -2614 474134
rect -2378 473898 586302 474134
rect 586538 473898 586622 474134
rect 586858 473898 592650 474134
rect -8726 473866 592650 473898
rect -8726 468174 592650 468206
rect -8726 467938 -1974 468174
rect -1738 467938 -1654 468174
rect -1418 467938 585342 468174
rect 585578 467938 585662 468174
rect 585898 467938 592650 468174
rect -8726 467854 592650 467938
rect -8726 467618 -1974 467854
rect -1738 467618 -1654 467854
rect -1418 467618 585342 467854
rect 585578 467618 585662 467854
rect 585898 467618 592650 467854
rect -8726 467586 592650 467618
rect -8726 464454 592650 464486
rect -8726 464218 -2934 464454
rect -2698 464218 -2614 464454
rect -2378 464218 586302 464454
rect 586538 464218 586622 464454
rect 586858 464218 592650 464454
rect -8726 464134 592650 464218
rect -8726 463898 -2934 464134
rect -2698 463898 -2614 464134
rect -2378 463898 586302 464134
rect 586538 463898 586622 464134
rect 586858 463898 592650 464134
rect -8726 463866 592650 463898
rect -8726 458174 592650 458206
rect -8726 457938 -1974 458174
rect -1738 457938 -1654 458174
rect -1418 457938 585342 458174
rect 585578 457938 585662 458174
rect 585898 457938 592650 458174
rect -8726 457854 592650 457938
rect -8726 457618 -1974 457854
rect -1738 457618 -1654 457854
rect -1418 457618 585342 457854
rect 585578 457618 585662 457854
rect 585898 457618 592650 457854
rect -8726 457586 592650 457618
rect -8726 454454 592650 454486
rect -8726 454218 -2934 454454
rect -2698 454218 -2614 454454
rect -2378 454218 586302 454454
rect 586538 454218 586622 454454
rect 586858 454218 592650 454454
rect -8726 454134 592650 454218
rect -8726 453898 -2934 454134
rect -2698 453898 -2614 454134
rect -2378 453898 586302 454134
rect 586538 453898 586622 454134
rect 586858 453898 592650 454134
rect -8726 453866 592650 453898
rect -8726 448174 592650 448206
rect -8726 447938 -1974 448174
rect -1738 447938 -1654 448174
rect -1418 447938 585342 448174
rect 585578 447938 585662 448174
rect 585898 447938 592650 448174
rect -8726 447854 592650 447938
rect -8726 447618 -1974 447854
rect -1738 447618 -1654 447854
rect -1418 447618 585342 447854
rect 585578 447618 585662 447854
rect 585898 447618 592650 447854
rect -8726 447586 592650 447618
rect -8726 444454 592650 444486
rect -8726 444218 -2934 444454
rect -2698 444218 -2614 444454
rect -2378 444218 586302 444454
rect 586538 444218 586622 444454
rect 586858 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -2934 444134
rect -2698 443898 -2614 444134
rect -2378 443898 586302 444134
rect 586538 443898 586622 444134
rect 586858 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 438174 592650 438206
rect -8726 437938 -1974 438174
rect -1738 437938 -1654 438174
rect -1418 437938 585342 438174
rect 585578 437938 585662 438174
rect 585898 437938 592650 438174
rect -8726 437854 592650 437938
rect -8726 437618 -1974 437854
rect -1738 437618 -1654 437854
rect -1418 437618 585342 437854
rect 585578 437618 585662 437854
rect 585898 437618 592650 437854
rect -8726 437586 592650 437618
rect -8726 434454 592650 434486
rect -8726 434218 -2934 434454
rect -2698 434218 -2614 434454
rect -2378 434218 586302 434454
rect 586538 434218 586622 434454
rect 586858 434218 592650 434454
rect -8726 434134 592650 434218
rect -8726 433898 -2934 434134
rect -2698 433898 -2614 434134
rect -2378 433898 586302 434134
rect 586538 433898 586622 434134
rect 586858 433898 592650 434134
rect -8726 433866 592650 433898
rect -8726 428174 592650 428206
rect -8726 427938 -1974 428174
rect -1738 427938 -1654 428174
rect -1418 427938 585342 428174
rect 585578 427938 585662 428174
rect 585898 427938 592650 428174
rect -8726 427854 592650 427938
rect -8726 427618 -1974 427854
rect -1738 427618 -1654 427854
rect -1418 427618 585342 427854
rect 585578 427618 585662 427854
rect 585898 427618 592650 427854
rect -8726 427586 592650 427618
rect -8726 424454 592650 424486
rect -8726 424218 -2934 424454
rect -2698 424218 -2614 424454
rect -2378 424218 586302 424454
rect 586538 424218 586622 424454
rect 586858 424218 592650 424454
rect -8726 424134 592650 424218
rect -8726 423898 -2934 424134
rect -2698 423898 -2614 424134
rect -2378 423898 586302 424134
rect 586538 423898 586622 424134
rect 586858 423898 592650 424134
rect -8726 423866 592650 423898
rect -8726 418174 592650 418206
rect -8726 417938 -1974 418174
rect -1738 417938 -1654 418174
rect -1418 417938 585342 418174
rect 585578 417938 585662 418174
rect 585898 417938 592650 418174
rect -8726 417854 592650 417938
rect -8726 417618 -1974 417854
rect -1738 417618 -1654 417854
rect -1418 417618 585342 417854
rect 585578 417618 585662 417854
rect 585898 417618 592650 417854
rect -8726 417586 592650 417618
rect -8726 414454 592650 414486
rect -8726 414218 -2934 414454
rect -2698 414218 -2614 414454
rect -2378 414218 586302 414454
rect 586538 414218 586622 414454
rect 586858 414218 592650 414454
rect -8726 414134 592650 414218
rect -8726 413898 -2934 414134
rect -2698 413898 -2614 414134
rect -2378 413898 586302 414134
rect 586538 413898 586622 414134
rect 586858 413898 592650 414134
rect -8726 413866 592650 413898
rect -8726 408174 592650 408206
rect -8726 407938 -1974 408174
rect -1738 407938 -1654 408174
rect -1418 407938 585342 408174
rect 585578 407938 585662 408174
rect 585898 407938 592650 408174
rect -8726 407854 592650 407938
rect -8726 407618 -1974 407854
rect -1738 407618 -1654 407854
rect -1418 407618 585342 407854
rect 585578 407618 585662 407854
rect 585898 407618 592650 407854
rect -8726 407586 592650 407618
rect -8726 404454 592650 404486
rect -8726 404218 -2934 404454
rect -2698 404218 -2614 404454
rect -2378 404218 586302 404454
rect 586538 404218 586622 404454
rect 586858 404218 592650 404454
rect -8726 404134 592650 404218
rect -8726 403898 -2934 404134
rect -2698 403898 -2614 404134
rect -2378 403898 586302 404134
rect 586538 403898 586622 404134
rect 586858 403898 592650 404134
rect -8726 403866 592650 403898
rect -8726 398174 592650 398206
rect -8726 397938 -1974 398174
rect -1738 397938 -1654 398174
rect -1418 397938 585342 398174
rect 585578 397938 585662 398174
rect 585898 397938 592650 398174
rect -8726 397854 592650 397938
rect -8726 397618 -1974 397854
rect -1738 397618 -1654 397854
rect -1418 397618 585342 397854
rect 585578 397618 585662 397854
rect 585898 397618 592650 397854
rect -8726 397586 592650 397618
rect -8726 394454 592650 394486
rect -8726 394218 -2934 394454
rect -2698 394218 -2614 394454
rect -2378 394218 586302 394454
rect 586538 394218 586622 394454
rect 586858 394218 592650 394454
rect -8726 394134 592650 394218
rect -8726 393898 -2934 394134
rect -2698 393898 -2614 394134
rect -2378 393898 586302 394134
rect 586538 393898 586622 394134
rect 586858 393898 592650 394134
rect -8726 393866 592650 393898
rect -8726 388174 592650 388206
rect -8726 387938 -1974 388174
rect -1738 387938 -1654 388174
rect -1418 387938 585342 388174
rect 585578 387938 585662 388174
rect 585898 387938 592650 388174
rect -8726 387854 592650 387938
rect -8726 387618 -1974 387854
rect -1738 387618 -1654 387854
rect -1418 387618 585342 387854
rect 585578 387618 585662 387854
rect 585898 387618 592650 387854
rect -8726 387586 592650 387618
rect -8726 384454 592650 384486
rect -8726 384218 -2934 384454
rect -2698 384218 -2614 384454
rect -2378 384218 586302 384454
rect 586538 384218 586622 384454
rect 586858 384218 592650 384454
rect -8726 384134 592650 384218
rect -8726 383898 -2934 384134
rect -2698 383898 -2614 384134
rect -2378 383898 586302 384134
rect 586538 383898 586622 384134
rect 586858 383898 592650 384134
rect -8726 383866 592650 383898
rect -8726 378174 592650 378206
rect -8726 377938 -1974 378174
rect -1738 377938 -1654 378174
rect -1418 377938 585342 378174
rect 585578 377938 585662 378174
rect 585898 377938 592650 378174
rect -8726 377854 592650 377938
rect -8726 377618 -1974 377854
rect -1738 377618 -1654 377854
rect -1418 377618 585342 377854
rect 585578 377618 585662 377854
rect 585898 377618 592650 377854
rect -8726 377586 592650 377618
rect -8726 374454 592650 374486
rect -8726 374218 -2934 374454
rect -2698 374218 -2614 374454
rect -2378 374218 586302 374454
rect 586538 374218 586622 374454
rect 586858 374218 592650 374454
rect -8726 374134 592650 374218
rect -8726 373898 -2934 374134
rect -2698 373898 -2614 374134
rect -2378 373898 586302 374134
rect 586538 373898 586622 374134
rect 586858 373898 592650 374134
rect -8726 373866 592650 373898
rect -8726 368174 592650 368206
rect -8726 367938 -1974 368174
rect -1738 367938 -1654 368174
rect -1418 367938 585342 368174
rect 585578 367938 585662 368174
rect 585898 367938 592650 368174
rect -8726 367854 592650 367938
rect -8726 367618 -1974 367854
rect -1738 367618 -1654 367854
rect -1418 367618 585342 367854
rect 585578 367618 585662 367854
rect 585898 367618 592650 367854
rect -8726 367586 592650 367618
rect -8726 364454 592650 364486
rect -8726 364218 -2934 364454
rect -2698 364218 -2614 364454
rect -2378 364218 586302 364454
rect 586538 364218 586622 364454
rect 586858 364218 592650 364454
rect -8726 364134 592650 364218
rect -8726 363898 -2934 364134
rect -2698 363898 -2614 364134
rect -2378 363898 586302 364134
rect 586538 363898 586622 364134
rect 586858 363898 592650 364134
rect -8726 363866 592650 363898
rect -8726 358174 592650 358206
rect -8726 357938 -1974 358174
rect -1738 357938 -1654 358174
rect -1418 357938 585342 358174
rect 585578 357938 585662 358174
rect 585898 357938 592650 358174
rect -8726 357854 592650 357938
rect -8726 357618 -1974 357854
rect -1738 357618 -1654 357854
rect -1418 357618 585342 357854
rect 585578 357618 585662 357854
rect 585898 357618 592650 357854
rect -8726 357586 592650 357618
rect -8726 354454 592650 354486
rect -8726 354218 -2934 354454
rect -2698 354218 -2614 354454
rect -2378 354218 586302 354454
rect 586538 354218 586622 354454
rect 586858 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -2934 354134
rect -2698 353898 -2614 354134
rect -2378 353898 586302 354134
rect 586538 353898 586622 354134
rect 586858 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 348174 592650 348206
rect -8726 347938 -1974 348174
rect -1738 347938 -1654 348174
rect -1418 347938 585342 348174
rect 585578 347938 585662 348174
rect 585898 347938 592650 348174
rect -8726 347854 592650 347938
rect -8726 347618 -1974 347854
rect -1738 347618 -1654 347854
rect -1418 347618 585342 347854
rect 585578 347618 585662 347854
rect 585898 347618 592650 347854
rect -8726 347586 592650 347618
rect -8726 344454 592650 344486
rect -8726 344218 -2934 344454
rect -2698 344218 -2614 344454
rect -2378 344218 586302 344454
rect 586538 344218 586622 344454
rect 586858 344218 592650 344454
rect -8726 344134 592650 344218
rect -8726 343898 -2934 344134
rect -2698 343898 -2614 344134
rect -2378 343898 586302 344134
rect 586538 343898 586622 344134
rect 586858 343898 592650 344134
rect -8726 343866 592650 343898
rect -8726 338174 592650 338206
rect -8726 337938 -1974 338174
rect -1738 337938 -1654 338174
rect -1418 337938 585342 338174
rect 585578 337938 585662 338174
rect 585898 337938 592650 338174
rect -8726 337854 592650 337938
rect -8726 337618 -1974 337854
rect -1738 337618 -1654 337854
rect -1418 337618 585342 337854
rect 585578 337618 585662 337854
rect 585898 337618 592650 337854
rect -8726 337586 592650 337618
rect -8726 334454 592650 334486
rect -8726 334218 -2934 334454
rect -2698 334218 -2614 334454
rect -2378 334218 586302 334454
rect 586538 334218 586622 334454
rect 586858 334218 592650 334454
rect -8726 334134 592650 334218
rect -8726 333898 -2934 334134
rect -2698 333898 -2614 334134
rect -2378 333898 586302 334134
rect 586538 333898 586622 334134
rect 586858 333898 592650 334134
rect -8726 333866 592650 333898
rect -8726 328174 592650 328206
rect -8726 327938 -1974 328174
rect -1738 327938 -1654 328174
rect -1418 327938 585342 328174
rect 585578 327938 585662 328174
rect 585898 327938 592650 328174
rect -8726 327854 592650 327938
rect -8726 327618 -1974 327854
rect -1738 327618 -1654 327854
rect -1418 327618 585342 327854
rect 585578 327618 585662 327854
rect 585898 327618 592650 327854
rect -8726 327586 592650 327618
rect -8726 324454 592650 324486
rect -8726 324218 -2934 324454
rect -2698 324218 -2614 324454
rect -2378 324218 586302 324454
rect 586538 324218 586622 324454
rect 586858 324218 592650 324454
rect -8726 324134 592650 324218
rect -8726 323898 -2934 324134
rect -2698 323898 -2614 324134
rect -2378 323898 586302 324134
rect 586538 323898 586622 324134
rect 586858 323898 592650 324134
rect -8726 323866 592650 323898
rect -8726 318174 592650 318206
rect -8726 317938 -1974 318174
rect -1738 317938 -1654 318174
rect -1418 317938 303504 318174
rect 303740 317938 437872 318174
rect 438108 317938 585342 318174
rect 585578 317938 585662 318174
rect 585898 317938 592650 318174
rect -8726 317854 592650 317938
rect -8726 317618 -1974 317854
rect -1738 317618 -1654 317854
rect -1418 317618 303504 317854
rect 303740 317618 437872 317854
rect 438108 317618 585342 317854
rect 585578 317618 585662 317854
rect 585898 317618 592650 317854
rect -8726 317586 592650 317618
rect -8726 314454 592650 314486
rect -8726 314218 -2934 314454
rect -2698 314218 -2614 314454
rect -2378 314218 302824 314454
rect 303060 314218 438552 314454
rect 438788 314218 586302 314454
rect 586538 314218 586622 314454
rect 586858 314218 592650 314454
rect -8726 314134 592650 314218
rect -8726 313898 -2934 314134
rect -2698 313898 -2614 314134
rect -2378 313898 302824 314134
rect 303060 313898 438552 314134
rect 438788 313898 586302 314134
rect 586538 313898 586622 314134
rect 586858 313898 592650 314134
rect -8726 313866 592650 313898
rect -8726 308174 592650 308206
rect -8726 307938 -1974 308174
rect -1738 307938 -1654 308174
rect -1418 307938 303504 308174
rect 303740 307938 437872 308174
rect 438108 307938 585342 308174
rect 585578 307938 585662 308174
rect 585898 307938 592650 308174
rect -8726 307854 592650 307938
rect -8726 307618 -1974 307854
rect -1738 307618 -1654 307854
rect -1418 307618 303504 307854
rect 303740 307618 437872 307854
rect 438108 307618 585342 307854
rect 585578 307618 585662 307854
rect 585898 307618 592650 307854
rect -8726 307586 592650 307618
rect -8726 304454 592650 304486
rect -8726 304218 -2934 304454
rect -2698 304218 -2614 304454
rect -2378 304218 302824 304454
rect 303060 304218 438552 304454
rect 438788 304218 586302 304454
rect 586538 304218 586622 304454
rect 586858 304218 592650 304454
rect -8726 304134 592650 304218
rect -8726 303898 -2934 304134
rect -2698 303898 -2614 304134
rect -2378 303898 302824 304134
rect 303060 303898 438552 304134
rect 438788 303898 586302 304134
rect 586538 303898 586622 304134
rect 586858 303898 592650 304134
rect -8726 303866 592650 303898
rect -8726 298174 592650 298206
rect -8726 297938 -1974 298174
rect -1738 297938 -1654 298174
rect -1418 297938 303504 298174
rect 303740 297938 437872 298174
rect 438108 297938 585342 298174
rect 585578 297938 585662 298174
rect 585898 297938 592650 298174
rect -8726 297854 592650 297938
rect -8726 297618 -1974 297854
rect -1738 297618 -1654 297854
rect -1418 297618 303504 297854
rect 303740 297618 437872 297854
rect 438108 297618 585342 297854
rect 585578 297618 585662 297854
rect 585898 297618 592650 297854
rect -8726 297586 592650 297618
rect -8726 294454 592650 294486
rect -8726 294218 -2934 294454
rect -2698 294218 -2614 294454
rect -2378 294218 302824 294454
rect 303060 294218 438552 294454
rect 438788 294218 586302 294454
rect 586538 294218 586622 294454
rect 586858 294218 592650 294454
rect -8726 294134 592650 294218
rect -8726 293898 -2934 294134
rect -2698 293898 -2614 294134
rect -2378 293898 302824 294134
rect 303060 293898 438552 294134
rect 438788 293898 586302 294134
rect 586538 293898 586622 294134
rect 586858 293898 592650 294134
rect -8726 293866 592650 293898
rect -8726 288174 592650 288206
rect -8726 287938 -1974 288174
rect -1738 287938 -1654 288174
rect -1418 287938 303504 288174
rect 303740 287938 437872 288174
rect 438108 287938 585342 288174
rect 585578 287938 585662 288174
rect 585898 287938 592650 288174
rect -8726 287854 592650 287938
rect -8726 287618 -1974 287854
rect -1738 287618 -1654 287854
rect -1418 287618 303504 287854
rect 303740 287618 437872 287854
rect 438108 287618 585342 287854
rect 585578 287618 585662 287854
rect 585898 287618 592650 287854
rect -8726 287586 592650 287618
rect -8726 284454 592650 284486
rect -8726 284218 -2934 284454
rect -2698 284218 -2614 284454
rect -2378 284218 302824 284454
rect 303060 284218 438552 284454
rect 438788 284218 586302 284454
rect 586538 284218 586622 284454
rect 586858 284218 592650 284454
rect -8726 284134 592650 284218
rect -8726 283898 -2934 284134
rect -2698 283898 -2614 284134
rect -2378 283898 302824 284134
rect 303060 283898 438552 284134
rect 438788 283898 586302 284134
rect 586538 283898 586622 284134
rect 586858 283898 592650 284134
rect -8726 283866 592650 283898
rect -8726 278174 592650 278206
rect -8726 277938 -1974 278174
rect -1738 277938 -1654 278174
rect -1418 277938 303504 278174
rect 303740 277938 437872 278174
rect 438108 277938 585342 278174
rect 585578 277938 585662 278174
rect 585898 277938 592650 278174
rect -8726 277927 592650 277938
rect -8726 277854 81714 277927
rect -8726 277618 -1974 277854
rect -1738 277618 -1654 277854
rect -1418 277691 81714 277854
rect 81950 277691 112434 277927
rect 112670 277691 143154 277927
rect 143390 277691 149978 277927
rect 150214 277691 180698 277927
rect 180934 277691 211418 277927
rect 211654 277854 592650 277927
rect 211654 277691 303504 277854
rect -1418 277618 303504 277691
rect 303740 277618 437872 277854
rect 438108 277618 585342 277854
rect 585578 277618 585662 277854
rect 585898 277618 592650 277854
rect -8726 277586 592650 277618
rect -8726 274454 592650 274486
rect -8726 274218 -2934 274454
rect -2698 274218 -2614 274454
rect -2378 274218 97074 274454
rect 97310 274218 127794 274454
rect 128030 274218 165338 274454
rect 165574 274218 196058 274454
rect 196294 274218 302824 274454
rect 303060 274218 438552 274454
rect 438788 274218 586302 274454
rect 586538 274218 586622 274454
rect 586858 274218 592650 274454
rect -8726 274134 592650 274218
rect -8726 273898 -2934 274134
rect -2698 273898 -2614 274134
rect -2378 273898 97074 274134
rect 97310 273898 127794 274134
rect 128030 273898 165338 274134
rect 165574 273898 196058 274134
rect 196294 273898 302824 274134
rect 303060 273898 438552 274134
rect 438788 273898 586302 274134
rect 586538 273898 586622 274134
rect 586858 273898 592650 274134
rect -8726 273866 592650 273898
rect -8726 268174 592650 268206
rect -8726 267938 -1974 268174
rect -1738 267938 -1654 268174
rect -1418 267938 81714 268174
rect 81950 267938 112434 268174
rect 112670 267938 143154 268174
rect 143390 267938 149978 268174
rect 150214 267938 180698 268174
rect 180934 267938 211418 268174
rect 211654 267938 303504 268174
rect 303740 267938 437872 268174
rect 438108 267938 585342 268174
rect 585578 267938 585662 268174
rect 585898 267938 592650 268174
rect -8726 267854 592650 267938
rect -8726 267618 -1974 267854
rect -1738 267618 -1654 267854
rect -1418 267618 81714 267854
rect 81950 267618 112434 267854
rect 112670 267618 143154 267854
rect 143390 267618 149978 267854
rect 150214 267618 180698 267854
rect 180934 267618 211418 267854
rect 211654 267618 303504 267854
rect 303740 267618 437872 267854
rect 438108 267618 585342 267854
rect 585578 267618 585662 267854
rect 585898 267618 592650 267854
rect -8726 267586 592650 267618
rect -8726 264454 592650 264486
rect -8726 264218 -2934 264454
rect -2698 264218 -2614 264454
rect -2378 264218 97074 264454
rect 97310 264218 127794 264454
rect 128030 264218 165338 264454
rect 165574 264218 196058 264454
rect 196294 264218 302824 264454
rect 303060 264218 438552 264454
rect 438788 264218 586302 264454
rect 586538 264218 586622 264454
rect 586858 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -2934 264134
rect -2698 263898 -2614 264134
rect -2378 263898 97074 264134
rect 97310 263898 127794 264134
rect 128030 263898 165338 264134
rect 165574 263898 196058 264134
rect 196294 263898 302824 264134
rect 303060 263898 438552 264134
rect 438788 263898 586302 264134
rect 586538 263898 586622 264134
rect 586858 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 258174 592650 258206
rect -8726 257938 -1974 258174
rect -1738 257938 -1654 258174
rect -1418 257938 81714 258174
rect 81950 257938 112434 258174
rect 112670 257938 143154 258174
rect 143390 257938 149978 258174
rect 150214 257938 180698 258174
rect 180934 257938 211418 258174
rect 211654 257938 303504 258174
rect 303740 257938 437872 258174
rect 438108 257938 585342 258174
rect 585578 257938 585662 258174
rect 585898 257938 592650 258174
rect -8726 257854 592650 257938
rect -8726 257618 -1974 257854
rect -1738 257618 -1654 257854
rect -1418 257618 81714 257854
rect 81950 257618 112434 257854
rect 112670 257618 143154 257854
rect 143390 257618 149978 257854
rect 150214 257618 180698 257854
rect 180934 257618 211418 257854
rect 211654 257618 303504 257854
rect 303740 257618 437872 257854
rect 438108 257618 585342 257854
rect 585578 257618 585662 257854
rect 585898 257618 592650 257854
rect -8726 257586 592650 257618
rect -8726 254454 592650 254486
rect -8726 254218 -2934 254454
rect -2698 254218 -2614 254454
rect -2378 254218 97074 254454
rect 97310 254218 127794 254454
rect 128030 254218 165338 254454
rect 165574 254218 196058 254454
rect 196294 254218 302824 254454
rect 303060 254218 438552 254454
rect 438788 254218 586302 254454
rect 586538 254218 586622 254454
rect 586858 254218 592650 254454
rect -8726 254134 592650 254218
rect -8726 253898 -2934 254134
rect -2698 253898 -2614 254134
rect -2378 253898 97074 254134
rect 97310 253898 127794 254134
rect 128030 253898 165338 254134
rect 165574 253898 196058 254134
rect 196294 253898 302824 254134
rect 303060 253898 438552 254134
rect 438788 253898 586302 254134
rect 586538 253898 586622 254134
rect 586858 253898 592650 254134
rect -8726 253866 592650 253898
rect -8726 248174 592650 248206
rect -8726 247938 -1974 248174
rect -1738 247938 -1654 248174
rect -1418 247938 81714 248174
rect 81950 247938 112434 248174
rect 112670 247938 143154 248174
rect 143390 247938 149978 248174
rect 150214 247938 180698 248174
rect 180934 247938 211418 248174
rect 211654 247938 303504 248174
rect 303740 247938 437872 248174
rect 438108 247938 585342 248174
rect 585578 247938 585662 248174
rect 585898 247938 592650 248174
rect -8726 247854 592650 247938
rect -8726 247618 -1974 247854
rect -1738 247618 -1654 247854
rect -1418 247618 81714 247854
rect 81950 247618 112434 247854
rect 112670 247618 143154 247854
rect 143390 247618 149978 247854
rect 150214 247618 180698 247854
rect 180934 247618 211418 247854
rect 211654 247618 303504 247854
rect 303740 247618 437872 247854
rect 438108 247618 585342 247854
rect 585578 247618 585662 247854
rect 585898 247618 592650 247854
rect -8726 247586 592650 247618
rect -8726 244454 592650 244486
rect -8726 244218 -2934 244454
rect -2698 244218 -2614 244454
rect -2378 244218 97074 244454
rect 97310 244218 127794 244454
rect 128030 244218 165338 244454
rect 165574 244218 196058 244454
rect 196294 244218 302824 244454
rect 303060 244218 438552 244454
rect 438788 244218 586302 244454
rect 586538 244218 586622 244454
rect 586858 244218 592650 244454
rect -8726 244134 592650 244218
rect -8726 243898 -2934 244134
rect -2698 243898 -2614 244134
rect -2378 243898 97074 244134
rect 97310 243898 127794 244134
rect 128030 243898 165338 244134
rect 165574 243898 196058 244134
rect 196294 243898 302824 244134
rect 303060 243898 438552 244134
rect 438788 243898 586302 244134
rect 586538 243898 586622 244134
rect 586858 243898 592650 244134
rect -8726 243866 592650 243898
rect -8726 238174 592650 238206
rect -8726 237938 -1974 238174
rect -1738 237938 -1654 238174
rect -1418 237938 81714 238174
rect 81950 237938 112434 238174
rect 112670 237938 143154 238174
rect 143390 237938 149978 238174
rect 150214 237938 180698 238174
rect 180934 237938 211418 238174
rect 211654 237938 585342 238174
rect 585578 237938 585662 238174
rect 585898 237938 592650 238174
rect -8726 237854 592650 237938
rect -8726 237618 -1974 237854
rect -1738 237618 -1654 237854
rect -1418 237618 81714 237854
rect 81950 237618 112434 237854
rect 112670 237618 143154 237854
rect 143390 237618 149978 237854
rect 150214 237618 180698 237854
rect 180934 237618 211418 237854
rect 211654 237618 585342 237854
rect 585578 237618 585662 237854
rect 585898 237618 592650 237854
rect -8726 237586 592650 237618
rect -8726 234454 592650 234486
rect -8726 234218 -2934 234454
rect -2698 234218 -2614 234454
rect -2378 234218 586302 234454
rect 586538 234218 586622 234454
rect 586858 234218 592650 234454
rect -8726 234134 592650 234218
rect -8726 233898 -2934 234134
rect -2698 233898 -2614 234134
rect -2378 233898 586302 234134
rect 586538 233898 586622 234134
rect 586858 233898 592650 234134
rect -8726 233866 592650 233898
rect -8726 228174 592650 228206
rect -8726 227938 -1974 228174
rect -1738 227938 -1654 228174
rect -1418 227938 116503 228174
rect 116739 227938 124345 228174
rect 124581 227938 132187 228174
rect 132423 227938 140029 228174
rect 140265 227938 409803 228174
rect 410039 227938 417645 228174
rect 417881 227938 425487 228174
rect 425723 227938 433329 228174
rect 433565 227938 585342 228174
rect 585578 227938 585662 228174
rect 585898 227938 592650 228174
rect -8726 227854 592650 227938
rect -8726 227618 -1974 227854
rect -1738 227618 -1654 227854
rect -1418 227618 116503 227854
rect 116739 227618 124345 227854
rect 124581 227618 132187 227854
rect 132423 227618 140029 227854
rect 140265 227618 409803 227854
rect 410039 227618 417645 227854
rect 417881 227618 425487 227854
rect 425723 227618 433329 227854
rect 433565 227618 585342 227854
rect 585578 227618 585662 227854
rect 585898 227618 592650 227854
rect -8726 227586 592650 227618
rect -8726 224454 592650 224486
rect -8726 224218 -2934 224454
rect -2698 224218 -2614 224454
rect -2378 224218 120424 224454
rect 120660 224218 128266 224454
rect 128502 224218 136108 224454
rect 136344 224218 143950 224454
rect 144186 224218 405882 224454
rect 406118 224218 413724 224454
rect 413960 224218 421566 224454
rect 421802 224218 429408 224454
rect 429644 224218 586302 224454
rect 586538 224218 586622 224454
rect 586858 224218 592650 224454
rect -8726 224134 592650 224218
rect -8726 223898 -2934 224134
rect -2698 223898 -2614 224134
rect -2378 223898 120424 224134
rect 120660 223898 128266 224134
rect 128502 223898 136108 224134
rect 136344 223898 143950 224134
rect 144186 223898 405882 224134
rect 406118 223898 413724 224134
rect 413960 223898 421566 224134
rect 421802 223898 429408 224134
rect 429644 223898 586302 224134
rect 586538 223898 586622 224134
rect 586858 223898 592650 224134
rect -8726 223866 592650 223898
rect -8726 218174 592650 218206
rect -8726 217938 -1974 218174
rect -1738 217938 -1654 218174
rect -1418 217938 116503 218174
rect 116739 217938 124345 218174
rect 124581 217938 132187 218174
rect 132423 217938 140029 218174
rect 140265 217938 409803 218174
rect 410039 217938 417645 218174
rect 417881 217938 425487 218174
rect 425723 217938 433329 218174
rect 433565 217938 585342 218174
rect 585578 217938 585662 218174
rect 585898 217938 592650 218174
rect -8726 217854 592650 217938
rect -8726 217618 -1974 217854
rect -1738 217618 -1654 217854
rect -1418 217618 116503 217854
rect 116739 217618 124345 217854
rect 124581 217618 132187 217854
rect 132423 217618 140029 217854
rect 140265 217618 409803 217854
rect 410039 217618 417645 217854
rect 417881 217618 425487 217854
rect 425723 217618 433329 217854
rect 433565 217618 585342 217854
rect 585578 217618 585662 217854
rect 585898 217618 592650 217854
rect -8726 217586 592650 217618
rect -8726 214454 592650 214486
rect -8726 214218 -2934 214454
rect -2698 214218 -2614 214454
rect -2378 214218 120424 214454
rect 120660 214218 128266 214454
rect 128502 214218 136108 214454
rect 136344 214218 143950 214454
rect 144186 214218 405882 214454
rect 406118 214218 413724 214454
rect 413960 214218 421566 214454
rect 421802 214218 429408 214454
rect 429644 214218 586302 214454
rect 586538 214218 586622 214454
rect 586858 214218 592650 214454
rect -8726 214134 592650 214218
rect -8726 213898 -2934 214134
rect -2698 213898 -2614 214134
rect -2378 213898 120424 214134
rect 120660 213898 128266 214134
rect 128502 213898 136108 214134
rect 136344 213898 143950 214134
rect 144186 213898 405882 214134
rect 406118 213898 413724 214134
rect 413960 213898 421566 214134
rect 421802 213898 429408 214134
rect 429644 213898 586302 214134
rect 586538 213898 586622 214134
rect 586858 213898 592650 214134
rect -8726 213866 592650 213898
rect -8726 208174 592650 208206
rect -8726 207938 -1974 208174
rect -1738 207938 -1654 208174
rect -1418 207938 14107 208174
rect 14343 207938 21949 208174
rect 22185 207938 29791 208174
rect 30027 207938 37633 208174
rect 37869 207938 42310 208174
rect 42546 207938 42630 208174
rect 42866 207938 42950 208174
rect 43186 207938 116503 208174
rect 116739 207938 124345 208174
rect 124581 207938 132187 208174
rect 132423 207938 140029 208174
rect 140265 207938 184767 208174
rect 185003 207938 192609 208174
rect 192845 207938 200451 208174
rect 200687 207938 208293 208174
rect 208529 207938 218899 208174
rect 219135 207938 226741 208174
rect 226977 207938 234583 208174
rect 234819 207938 242425 208174
rect 242661 207938 253031 208174
rect 253267 207938 260873 208174
rect 261109 207938 268715 208174
rect 268951 207938 276557 208174
rect 276793 207938 307407 208174
rect 307643 207938 315249 208174
rect 315485 207938 323091 208174
rect 323327 207938 330933 208174
rect 331169 207938 341539 208174
rect 341775 207938 349381 208174
rect 349617 207938 357223 208174
rect 357459 207938 365065 208174
rect 365301 207938 375671 208174
rect 375907 207938 383513 208174
rect 383749 207938 391355 208174
rect 391591 207938 399197 208174
rect 399433 207938 409803 208174
rect 410039 207938 417645 208174
rect 417881 207938 425487 208174
rect 425723 207938 433329 208174
rect 433565 207938 443935 208174
rect 444171 207938 451777 208174
rect 452013 207938 459619 208174
rect 459855 207938 467461 208174
rect 467697 207938 478067 208174
rect 478303 207938 485909 208174
rect 486145 207938 493751 208174
rect 493987 207938 501593 208174
rect 501829 207938 512199 208174
rect 512435 207938 520041 208174
rect 520277 207938 527883 208174
rect 528119 207938 535725 208174
rect 535961 207938 546331 208174
rect 546567 207938 554173 208174
rect 554409 207938 562015 208174
rect 562251 207938 569857 208174
rect 570093 207938 585342 208174
rect 585578 207938 585662 208174
rect 585898 207938 592650 208174
rect -8726 207854 592650 207938
rect -8726 207618 -1974 207854
rect -1738 207618 -1654 207854
rect -1418 207618 14107 207854
rect 14343 207618 21949 207854
rect 22185 207618 29791 207854
rect 30027 207618 37633 207854
rect 37869 207618 42310 207854
rect 42546 207618 42630 207854
rect 42866 207618 42950 207854
rect 43186 207618 116503 207854
rect 116739 207618 124345 207854
rect 124581 207618 132187 207854
rect 132423 207618 140029 207854
rect 140265 207618 184767 207854
rect 185003 207618 192609 207854
rect 192845 207618 200451 207854
rect 200687 207618 208293 207854
rect 208529 207618 218899 207854
rect 219135 207618 226741 207854
rect 226977 207618 234583 207854
rect 234819 207618 242425 207854
rect 242661 207618 253031 207854
rect 253267 207618 260873 207854
rect 261109 207618 268715 207854
rect 268951 207618 276557 207854
rect 276793 207618 307407 207854
rect 307643 207618 315249 207854
rect 315485 207618 323091 207854
rect 323327 207618 330933 207854
rect 331169 207618 341539 207854
rect 341775 207618 349381 207854
rect 349617 207618 357223 207854
rect 357459 207618 365065 207854
rect 365301 207618 375671 207854
rect 375907 207618 383513 207854
rect 383749 207618 391355 207854
rect 391591 207618 399197 207854
rect 399433 207618 409803 207854
rect 410039 207618 417645 207854
rect 417881 207618 425487 207854
rect 425723 207618 433329 207854
rect 433565 207618 443935 207854
rect 444171 207618 451777 207854
rect 452013 207618 459619 207854
rect 459855 207618 467461 207854
rect 467697 207618 478067 207854
rect 478303 207618 485909 207854
rect 486145 207618 493751 207854
rect 493987 207618 501593 207854
rect 501829 207618 512199 207854
rect 512435 207618 520041 207854
rect 520277 207618 527883 207854
rect 528119 207618 535725 207854
rect 535961 207618 546331 207854
rect 546567 207618 554173 207854
rect 554409 207618 562015 207854
rect 562251 207618 569857 207854
rect 570093 207618 585342 207854
rect 585578 207618 585662 207854
rect 585898 207618 592650 207854
rect -8726 207586 592650 207618
rect -8726 204454 592650 204486
rect -8726 204218 -2934 204454
rect -2698 204218 -2614 204454
rect -2378 204218 18028 204454
rect 18264 204218 25870 204454
rect 26106 204218 33712 204454
rect 33948 204218 41554 204454
rect 41790 204218 52160 204454
rect 52396 204218 60002 204454
rect 60238 204218 67844 204454
rect 68080 204218 75686 204454
rect 75922 204218 120424 204454
rect 120660 204218 128266 204454
rect 128502 204218 136108 204454
rect 136344 204218 143950 204454
rect 144186 204218 188688 204454
rect 188924 204218 196530 204454
rect 196766 204218 204372 204454
rect 204608 204218 212214 204454
rect 212450 204218 222820 204454
rect 223056 204218 230662 204454
rect 230898 204218 238504 204454
rect 238740 204218 246346 204454
rect 246582 204218 256952 204454
rect 257188 204218 264794 204454
rect 265030 204218 272636 204454
rect 272872 204218 280478 204454
rect 280714 204218 303486 204454
rect 303722 204218 311328 204454
rect 311564 204218 319170 204454
rect 319406 204218 327012 204454
rect 327248 204218 337618 204454
rect 337854 204218 345460 204454
rect 345696 204218 353302 204454
rect 353538 204218 361144 204454
rect 361380 204218 371750 204454
rect 371986 204218 379592 204454
rect 379828 204218 387434 204454
rect 387670 204218 395276 204454
rect 395512 204218 405882 204454
rect 406118 204218 413724 204454
rect 413960 204218 421566 204454
rect 421802 204218 429408 204454
rect 429644 204218 440014 204454
rect 440250 204218 447856 204454
rect 448092 204218 455698 204454
rect 455934 204218 463540 204454
rect 463776 204218 474146 204454
rect 474382 204218 481988 204454
rect 482224 204218 489830 204454
rect 490066 204218 497672 204454
rect 497908 204218 508278 204454
rect 508514 204218 516120 204454
rect 516356 204218 523962 204454
rect 524198 204218 531804 204454
rect 532040 204218 542410 204454
rect 542646 204218 550252 204454
rect 550488 204218 558094 204454
rect 558330 204218 565936 204454
rect 566172 204218 586302 204454
rect 586538 204218 586622 204454
rect 586858 204218 592650 204454
rect -8726 204134 592650 204218
rect -8726 203898 -2934 204134
rect -2698 203898 -2614 204134
rect -2378 203898 18028 204134
rect 18264 203898 25870 204134
rect 26106 203898 33712 204134
rect 33948 203898 41554 204134
rect 41790 203898 52160 204134
rect 52396 203898 60002 204134
rect 60238 203898 67844 204134
rect 68080 203898 75686 204134
rect 75922 203898 120424 204134
rect 120660 203898 128266 204134
rect 128502 203898 136108 204134
rect 136344 203898 143950 204134
rect 144186 203898 188688 204134
rect 188924 203898 196530 204134
rect 196766 203898 204372 204134
rect 204608 203898 212214 204134
rect 212450 203898 222820 204134
rect 223056 203898 230662 204134
rect 230898 203898 238504 204134
rect 238740 203898 246346 204134
rect 246582 203898 256952 204134
rect 257188 203898 264794 204134
rect 265030 203898 272636 204134
rect 272872 203898 280478 204134
rect 280714 203898 303486 204134
rect 303722 203898 311328 204134
rect 311564 203898 319170 204134
rect 319406 203898 327012 204134
rect 327248 203898 337618 204134
rect 337854 203898 345460 204134
rect 345696 203898 353302 204134
rect 353538 203898 361144 204134
rect 361380 203898 371750 204134
rect 371986 203898 379592 204134
rect 379828 203898 387434 204134
rect 387670 203898 395276 204134
rect 395512 203898 405882 204134
rect 406118 203898 413724 204134
rect 413960 203898 421566 204134
rect 421802 203898 429408 204134
rect 429644 203898 440014 204134
rect 440250 203898 447856 204134
rect 448092 203898 455698 204134
rect 455934 203898 463540 204134
rect 463776 203898 474146 204134
rect 474382 203898 481988 204134
rect 482224 203898 489830 204134
rect 490066 203898 497672 204134
rect 497908 203898 508278 204134
rect 508514 203898 516120 204134
rect 516356 203898 523962 204134
rect 524198 203898 531804 204134
rect 532040 203898 542410 204134
rect 542646 203898 550252 204134
rect 550488 203898 558094 204134
rect 558330 203898 565936 204134
rect 566172 203898 586302 204134
rect 586538 203898 586622 204134
rect 586858 203898 592650 204134
rect -8726 203866 592650 203898
rect -8726 198174 592650 198206
rect -8726 197938 -1974 198174
rect -1738 197938 -1654 198174
rect -1418 197938 14107 198174
rect 14343 197938 21949 198174
rect 22185 197938 29791 198174
rect 30027 197938 37633 198174
rect 37869 197938 42310 198174
rect 42546 197938 42630 198174
rect 42866 197938 42950 198174
rect 43186 197938 116503 198174
rect 116739 197938 124345 198174
rect 124581 197938 132187 198174
rect 132423 197938 140029 198174
rect 140265 197938 184767 198174
rect 185003 197938 192609 198174
rect 192845 197938 200451 198174
rect 200687 197938 208293 198174
rect 208529 197938 218899 198174
rect 219135 197938 226741 198174
rect 226977 197938 234583 198174
rect 234819 197938 242425 198174
rect 242661 197938 253031 198174
rect 253267 197938 260873 198174
rect 261109 197938 268715 198174
rect 268951 197938 276557 198174
rect 276793 197938 307407 198174
rect 307643 197938 315249 198174
rect 315485 197938 323091 198174
rect 323327 197938 330933 198174
rect 331169 197938 341539 198174
rect 341775 197938 349381 198174
rect 349617 197938 357223 198174
rect 357459 197938 365065 198174
rect 365301 197938 375671 198174
rect 375907 197938 383513 198174
rect 383749 197938 391355 198174
rect 391591 197938 399197 198174
rect 399433 197938 409803 198174
rect 410039 197938 417645 198174
rect 417881 197938 425487 198174
rect 425723 197938 433329 198174
rect 433565 197938 443935 198174
rect 444171 197938 451777 198174
rect 452013 197938 459619 198174
rect 459855 197938 467461 198174
rect 467697 197938 478067 198174
rect 478303 197938 485909 198174
rect 486145 197938 493751 198174
rect 493987 197938 501593 198174
rect 501829 197938 512199 198174
rect 512435 197938 520041 198174
rect 520277 197938 527883 198174
rect 528119 197938 535725 198174
rect 535961 197938 546331 198174
rect 546567 197938 554173 198174
rect 554409 197938 562015 198174
rect 562251 197938 569857 198174
rect 570093 197938 585342 198174
rect 585578 197938 585662 198174
rect 585898 197938 592650 198174
rect -8726 197854 592650 197938
rect -8726 197618 -1974 197854
rect -1738 197618 -1654 197854
rect -1418 197618 14107 197854
rect 14343 197618 21949 197854
rect 22185 197618 29791 197854
rect 30027 197618 37633 197854
rect 37869 197618 42310 197854
rect 42546 197618 42630 197854
rect 42866 197618 42950 197854
rect 43186 197618 116503 197854
rect 116739 197618 124345 197854
rect 124581 197618 132187 197854
rect 132423 197618 140029 197854
rect 140265 197618 184767 197854
rect 185003 197618 192609 197854
rect 192845 197618 200451 197854
rect 200687 197618 208293 197854
rect 208529 197618 218899 197854
rect 219135 197618 226741 197854
rect 226977 197618 234583 197854
rect 234819 197618 242425 197854
rect 242661 197618 253031 197854
rect 253267 197618 260873 197854
rect 261109 197618 268715 197854
rect 268951 197618 276557 197854
rect 276793 197618 307407 197854
rect 307643 197618 315249 197854
rect 315485 197618 323091 197854
rect 323327 197618 330933 197854
rect 331169 197618 341539 197854
rect 341775 197618 349381 197854
rect 349617 197618 357223 197854
rect 357459 197618 365065 197854
rect 365301 197618 375671 197854
rect 375907 197618 383513 197854
rect 383749 197618 391355 197854
rect 391591 197618 399197 197854
rect 399433 197618 409803 197854
rect 410039 197618 417645 197854
rect 417881 197618 425487 197854
rect 425723 197618 433329 197854
rect 433565 197618 443935 197854
rect 444171 197618 451777 197854
rect 452013 197618 459619 197854
rect 459855 197618 467461 197854
rect 467697 197618 478067 197854
rect 478303 197618 485909 197854
rect 486145 197618 493751 197854
rect 493987 197618 501593 197854
rect 501829 197618 512199 197854
rect 512435 197618 520041 197854
rect 520277 197618 527883 197854
rect 528119 197618 535725 197854
rect 535961 197618 546331 197854
rect 546567 197618 554173 197854
rect 554409 197618 562015 197854
rect 562251 197618 569857 197854
rect 570093 197618 585342 197854
rect 585578 197618 585662 197854
rect 585898 197618 592650 197854
rect -8726 197586 592650 197618
rect -8726 194454 592650 194486
rect -8726 194218 -2934 194454
rect -2698 194218 -2614 194454
rect -2378 194218 18028 194454
rect 18264 194218 25870 194454
rect 26106 194218 33712 194454
rect 33948 194218 41554 194454
rect 41790 194218 52160 194454
rect 52396 194218 60002 194454
rect 60238 194218 67844 194454
rect 68080 194218 75686 194454
rect 75922 194218 120424 194454
rect 120660 194218 128266 194454
rect 128502 194218 136108 194454
rect 136344 194218 143950 194454
rect 144186 194218 188688 194454
rect 188924 194218 196530 194454
rect 196766 194218 204372 194454
rect 204608 194218 212214 194454
rect 212450 194218 222820 194454
rect 223056 194218 230662 194454
rect 230898 194218 238504 194454
rect 238740 194218 246346 194454
rect 246582 194218 256952 194454
rect 257188 194218 264794 194454
rect 265030 194218 272636 194454
rect 272872 194218 280478 194454
rect 280714 194218 303486 194454
rect 303722 194218 311328 194454
rect 311564 194218 319170 194454
rect 319406 194218 327012 194454
rect 327248 194218 337618 194454
rect 337854 194218 345460 194454
rect 345696 194218 353302 194454
rect 353538 194218 361144 194454
rect 361380 194218 371750 194454
rect 371986 194218 379592 194454
rect 379828 194218 387434 194454
rect 387670 194218 395276 194454
rect 395512 194218 405882 194454
rect 406118 194218 413724 194454
rect 413960 194218 421566 194454
rect 421802 194218 429408 194454
rect 429644 194218 440014 194454
rect 440250 194218 447856 194454
rect 448092 194218 455698 194454
rect 455934 194218 463540 194454
rect 463776 194218 474146 194454
rect 474382 194218 481988 194454
rect 482224 194218 489830 194454
rect 490066 194218 497672 194454
rect 497908 194218 508278 194454
rect 508514 194218 516120 194454
rect 516356 194218 523962 194454
rect 524198 194218 531804 194454
rect 532040 194218 542410 194454
rect 542646 194218 550252 194454
rect 550488 194218 558094 194454
rect 558330 194218 565936 194454
rect 566172 194218 586302 194454
rect 586538 194218 586622 194454
rect 586858 194218 592650 194454
rect -8726 194134 592650 194218
rect -8726 193898 -2934 194134
rect -2698 193898 -2614 194134
rect -2378 193898 18028 194134
rect 18264 193898 25870 194134
rect 26106 193898 33712 194134
rect 33948 193898 41554 194134
rect 41790 193898 52160 194134
rect 52396 193898 60002 194134
rect 60238 193898 67844 194134
rect 68080 193898 75686 194134
rect 75922 193898 120424 194134
rect 120660 193898 128266 194134
rect 128502 193898 136108 194134
rect 136344 193898 143950 194134
rect 144186 193898 188688 194134
rect 188924 193898 196530 194134
rect 196766 193898 204372 194134
rect 204608 193898 212214 194134
rect 212450 193898 222820 194134
rect 223056 193898 230662 194134
rect 230898 193898 238504 194134
rect 238740 193898 246346 194134
rect 246582 193898 256952 194134
rect 257188 193898 264794 194134
rect 265030 193898 272636 194134
rect 272872 193898 280478 194134
rect 280714 193898 303486 194134
rect 303722 193898 311328 194134
rect 311564 193898 319170 194134
rect 319406 193898 327012 194134
rect 327248 193898 337618 194134
rect 337854 193898 345460 194134
rect 345696 193898 353302 194134
rect 353538 193898 361144 194134
rect 361380 193898 371750 194134
rect 371986 193898 379592 194134
rect 379828 193898 387434 194134
rect 387670 193898 395276 194134
rect 395512 193898 405882 194134
rect 406118 193898 413724 194134
rect 413960 193898 421566 194134
rect 421802 193898 429408 194134
rect 429644 193898 440014 194134
rect 440250 193898 447856 194134
rect 448092 193898 455698 194134
rect 455934 193898 463540 194134
rect 463776 193898 474146 194134
rect 474382 193898 481988 194134
rect 482224 193898 489830 194134
rect 490066 193898 497672 194134
rect 497908 193898 508278 194134
rect 508514 193898 516120 194134
rect 516356 193898 523962 194134
rect 524198 193898 531804 194134
rect 532040 193898 542410 194134
rect 542646 193898 550252 194134
rect 550488 193898 558094 194134
rect 558330 193898 565936 194134
rect 566172 193898 586302 194134
rect 586538 193898 586622 194134
rect 586858 193898 592650 194134
rect -8726 193866 592650 193898
rect -8726 188174 592650 188206
rect -8726 187938 -1974 188174
rect -1738 187938 -1654 188174
rect -1418 187938 43984 188174
rect 44220 187938 111581 188174
rect 111817 187938 179178 188174
rect 179414 187938 246775 188174
rect 247011 187938 337189 188174
rect 337425 187938 404786 188174
rect 405022 187938 472383 188174
rect 472619 187938 539980 188174
rect 540216 187938 585342 188174
rect 585578 187938 585662 188174
rect 585898 187938 592650 188174
rect -8726 187854 592650 187938
rect -8726 187618 -1974 187854
rect -1738 187618 -1654 187854
rect -1418 187618 43984 187854
rect 44220 187618 111581 187854
rect 111817 187618 179178 187854
rect 179414 187618 246775 187854
rect 247011 187618 337189 187854
rect 337425 187618 404786 187854
rect 405022 187618 472383 187854
rect 472619 187618 539980 187854
rect 540216 187618 585342 187854
rect 585578 187618 585662 187854
rect 585898 187618 592650 187854
rect -8726 187586 592650 187618
rect -8726 184454 592650 184486
rect -8726 184218 -2934 184454
rect -2698 184218 -2614 184454
rect -2378 184218 77782 184454
rect 78018 184218 145379 184454
rect 145615 184218 212976 184454
rect 213212 184218 280573 184454
rect 280809 184218 303391 184454
rect 303627 184218 370988 184454
rect 371224 184218 438585 184454
rect 438821 184218 506182 184454
rect 506418 184218 586302 184454
rect 586538 184218 586622 184454
rect 586858 184218 592650 184454
rect -8726 184134 592650 184218
rect -8726 183898 -2934 184134
rect -2698 183898 -2614 184134
rect -2378 183898 77782 184134
rect 78018 183898 145379 184134
rect 145615 183898 212976 184134
rect 213212 183898 280573 184134
rect 280809 183898 303391 184134
rect 303627 183898 370988 184134
rect 371224 183898 438585 184134
rect 438821 183898 506182 184134
rect 506418 183898 586302 184134
rect 586538 183898 586622 184134
rect 586858 183898 592650 184134
rect -8726 183866 592650 183898
rect -8726 178174 592650 178206
rect -8726 177938 -1974 178174
rect -1738 177938 -1654 178174
rect -1418 177938 585342 178174
rect 585578 177938 585662 178174
rect 585898 177938 592650 178174
rect -8726 177879 592650 177938
rect -8726 177854 48239 177879
rect -8726 177618 -1974 177854
rect -1738 177618 -1654 177854
rect -1418 177643 48239 177854
rect 48475 177643 56081 177879
rect 56317 177643 63923 177879
rect 64159 177643 71765 177879
rect 72001 177643 82371 177879
rect 82607 177643 90213 177879
rect 90449 177643 98055 177879
rect 98291 177643 105897 177879
rect 106133 177643 116503 177879
rect 116739 177643 124345 177879
rect 124581 177643 132187 177879
rect 132423 177643 140029 177879
rect 140265 177643 149978 177879
rect 150214 177643 180698 177879
rect 180934 177643 211418 177879
rect 211654 177643 242138 177879
rect 242374 177643 272858 177879
rect 273094 177643 307407 177879
rect 307643 177643 315249 177879
rect 315485 177643 323091 177879
rect 323327 177643 330933 177879
rect 331169 177643 341539 177879
rect 341775 177643 349381 177879
rect 349617 177643 357223 177879
rect 357459 177643 365065 177879
rect 365301 177643 375671 177879
rect 375907 177643 383513 177879
rect 383749 177643 391355 177879
rect 391591 177643 399197 177879
rect 399433 177643 443935 177879
rect 444171 177643 451777 177879
rect 452013 177643 459619 177879
rect 459855 177643 467461 177879
rect 467697 177643 478067 177879
rect 478303 177643 485909 177879
rect 486145 177643 493751 177879
rect 493987 177643 501593 177879
rect 501829 177643 512199 177879
rect 512435 177643 520041 177879
rect 520277 177643 527883 177879
rect 528119 177643 535725 177879
rect 535961 177854 592650 177879
rect 535961 177643 585342 177854
rect -1418 177618 585342 177643
rect 585578 177618 585662 177854
rect 585898 177618 592650 177854
rect -8726 177586 592650 177618
rect -8726 174454 592650 174486
rect -8726 174218 -2934 174454
rect -2698 174218 -2614 174454
rect -2378 174218 52160 174454
rect 52396 174218 60002 174454
rect 60238 174218 67844 174454
rect 68080 174218 75686 174454
rect 75922 174218 86292 174454
rect 86528 174218 94134 174454
rect 94370 174218 101976 174454
rect 102212 174218 109818 174454
rect 110054 174218 120424 174454
rect 120660 174218 128266 174454
rect 128502 174218 136108 174454
rect 136344 174218 143950 174454
rect 144186 174218 165338 174454
rect 165574 174218 196058 174454
rect 196294 174218 226778 174454
rect 227014 174218 257498 174454
rect 257734 174218 303486 174454
rect 303722 174218 311328 174454
rect 311564 174218 319170 174454
rect 319406 174218 327012 174454
rect 327248 174218 337618 174454
rect 337854 174218 345460 174454
rect 345696 174218 353302 174454
rect 353538 174218 361144 174454
rect 361380 174218 371750 174454
rect 371986 174218 379592 174454
rect 379828 174218 387434 174454
rect 387670 174218 395276 174454
rect 395512 174218 440014 174454
rect 440250 174218 447856 174454
rect 448092 174218 455698 174454
rect 455934 174218 463540 174454
rect 463776 174218 474146 174454
rect 474382 174218 481988 174454
rect 482224 174218 489830 174454
rect 490066 174218 497672 174454
rect 497908 174218 508278 174454
rect 508514 174218 516120 174454
rect 516356 174218 523962 174454
rect 524198 174218 531804 174454
rect 532040 174218 586302 174454
rect 586538 174218 586622 174454
rect 586858 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -2934 174134
rect -2698 173898 -2614 174134
rect -2378 173898 52160 174134
rect 52396 173898 60002 174134
rect 60238 173898 67844 174134
rect 68080 173898 75686 174134
rect 75922 173898 86292 174134
rect 86528 173898 94134 174134
rect 94370 173898 101976 174134
rect 102212 173898 109818 174134
rect 110054 173898 120424 174134
rect 120660 173898 128266 174134
rect 128502 173898 136108 174134
rect 136344 173898 143950 174134
rect 144186 173898 165338 174134
rect 165574 173898 196058 174134
rect 196294 173898 226778 174134
rect 227014 173898 257498 174134
rect 257734 173898 303486 174134
rect 303722 173898 311328 174134
rect 311564 173898 319170 174134
rect 319406 173898 327012 174134
rect 327248 173898 337618 174134
rect 337854 173898 345460 174134
rect 345696 173898 353302 174134
rect 353538 173898 361144 174134
rect 361380 173898 371750 174134
rect 371986 173898 379592 174134
rect 379828 173898 387434 174134
rect 387670 173898 395276 174134
rect 395512 173898 440014 174134
rect 440250 173898 447856 174134
rect 448092 173898 455698 174134
rect 455934 173898 463540 174134
rect 463776 173898 474146 174134
rect 474382 173898 481988 174134
rect 482224 173898 489830 174134
rect 490066 173898 497672 174134
rect 497908 173898 508278 174134
rect 508514 173898 516120 174134
rect 516356 173898 523962 174134
rect 524198 173898 531804 174134
rect 532040 173898 586302 174134
rect 586538 173898 586622 174134
rect 586858 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 168174 592650 168206
rect -8726 167938 -1974 168174
rect -1738 167938 -1654 168174
rect -1418 167938 48239 168174
rect 48475 167938 56081 168174
rect 56317 167938 63923 168174
rect 64159 167938 71765 168174
rect 72001 167938 82371 168174
rect 82607 167938 90213 168174
rect 90449 167938 98055 168174
rect 98291 167938 105897 168174
rect 106133 167938 116503 168174
rect 116739 167938 124345 168174
rect 124581 167938 132187 168174
rect 132423 167938 140029 168174
rect 140265 167938 149978 168174
rect 150214 167938 180698 168174
rect 180934 167938 211418 168174
rect 211654 167938 242138 168174
rect 242374 167938 272858 168174
rect 273094 167938 307407 168174
rect 307643 167938 315249 168174
rect 315485 167938 323091 168174
rect 323327 167938 330933 168174
rect 331169 167938 341539 168174
rect 341775 167938 349381 168174
rect 349617 167938 357223 168174
rect 357459 167938 365065 168174
rect 365301 167938 375671 168174
rect 375907 167938 383513 168174
rect 383749 167938 391355 168174
rect 391591 167938 399197 168174
rect 399433 167938 443935 168174
rect 444171 167938 451777 168174
rect 452013 167938 459619 168174
rect 459855 167938 467461 168174
rect 467697 167938 478067 168174
rect 478303 167938 485909 168174
rect 486145 167938 493751 168174
rect 493987 167938 501593 168174
rect 501829 167938 512199 168174
rect 512435 167938 520041 168174
rect 520277 167938 527883 168174
rect 528119 167938 535725 168174
rect 535961 167938 585342 168174
rect 585578 167938 585662 168174
rect 585898 167938 592650 168174
rect -8726 167854 592650 167938
rect -8726 167618 -1974 167854
rect -1738 167618 -1654 167854
rect -1418 167618 48239 167854
rect 48475 167618 56081 167854
rect 56317 167618 63923 167854
rect 64159 167618 71765 167854
rect 72001 167618 82371 167854
rect 82607 167618 90213 167854
rect 90449 167618 98055 167854
rect 98291 167618 105897 167854
rect 106133 167618 116503 167854
rect 116739 167618 124345 167854
rect 124581 167618 132187 167854
rect 132423 167618 140029 167854
rect 140265 167618 149978 167854
rect 150214 167618 180698 167854
rect 180934 167618 211418 167854
rect 211654 167618 242138 167854
rect 242374 167618 272858 167854
rect 273094 167618 307407 167854
rect 307643 167618 315249 167854
rect 315485 167618 323091 167854
rect 323327 167618 330933 167854
rect 331169 167618 341539 167854
rect 341775 167618 349381 167854
rect 349617 167618 357223 167854
rect 357459 167618 365065 167854
rect 365301 167618 375671 167854
rect 375907 167618 383513 167854
rect 383749 167618 391355 167854
rect 391591 167618 399197 167854
rect 399433 167618 443935 167854
rect 444171 167618 451777 167854
rect 452013 167618 459619 167854
rect 459855 167618 467461 167854
rect 467697 167618 478067 167854
rect 478303 167618 485909 167854
rect 486145 167618 493751 167854
rect 493987 167618 501593 167854
rect 501829 167618 512199 167854
rect 512435 167618 520041 167854
rect 520277 167618 527883 167854
rect 528119 167618 535725 167854
rect 535961 167618 585342 167854
rect 585578 167618 585662 167854
rect 585898 167618 592650 167854
rect -8726 167586 592650 167618
rect -8726 164454 592650 164486
rect -8726 164218 -2934 164454
rect -2698 164218 -2614 164454
rect -2378 164218 52160 164454
rect 52396 164218 60002 164454
rect 60238 164218 67844 164454
rect 68080 164218 75686 164454
rect 75922 164218 86292 164454
rect 86528 164218 94134 164454
rect 94370 164218 101976 164454
rect 102212 164218 109818 164454
rect 110054 164218 120424 164454
rect 120660 164218 128266 164454
rect 128502 164218 136108 164454
rect 136344 164218 143950 164454
rect 144186 164218 165338 164454
rect 165574 164218 196058 164454
rect 196294 164218 226778 164454
rect 227014 164218 257498 164454
rect 257734 164218 277814 164454
rect 278050 164218 303486 164454
rect 303722 164218 311328 164454
rect 311564 164218 319170 164454
rect 319406 164218 327012 164454
rect 327248 164218 337618 164454
rect 337854 164218 345460 164454
rect 345696 164218 353302 164454
rect 353538 164218 361144 164454
rect 361380 164218 371750 164454
rect 371986 164218 379592 164454
rect 379828 164218 387434 164454
rect 387670 164218 395276 164454
rect 395512 164218 440014 164454
rect 440250 164218 447856 164454
rect 448092 164218 455698 164454
rect 455934 164218 463540 164454
rect 463776 164218 474146 164454
rect 474382 164218 481988 164454
rect 482224 164218 489830 164454
rect 490066 164218 497672 164454
rect 497908 164218 508278 164454
rect 508514 164218 516120 164454
rect 516356 164218 523962 164454
rect 524198 164218 531804 164454
rect 532040 164218 586302 164454
rect 586538 164218 586622 164454
rect 586858 164218 592650 164454
rect -8726 164134 592650 164218
rect -8726 163898 -2934 164134
rect -2698 163898 -2614 164134
rect -2378 163898 52160 164134
rect 52396 163898 60002 164134
rect 60238 163898 67844 164134
rect 68080 163898 75686 164134
rect 75922 163898 86292 164134
rect 86528 163898 94134 164134
rect 94370 163898 101976 164134
rect 102212 163898 109818 164134
rect 110054 163898 120424 164134
rect 120660 163898 128266 164134
rect 128502 163898 136108 164134
rect 136344 163898 143950 164134
rect 144186 163898 165338 164134
rect 165574 163898 196058 164134
rect 196294 163898 226778 164134
rect 227014 163898 257498 164134
rect 257734 163898 277814 164134
rect 278050 163898 303486 164134
rect 303722 163898 311328 164134
rect 311564 163898 319170 164134
rect 319406 163898 327012 164134
rect 327248 163898 337618 164134
rect 337854 163898 345460 164134
rect 345696 163898 353302 164134
rect 353538 163898 361144 164134
rect 361380 163898 371750 164134
rect 371986 163898 379592 164134
rect 379828 163898 387434 164134
rect 387670 163898 395276 164134
rect 395512 163898 440014 164134
rect 440250 163898 447856 164134
rect 448092 163898 455698 164134
rect 455934 163898 463540 164134
rect 463776 163898 474146 164134
rect 474382 163898 481988 164134
rect 482224 163898 489830 164134
rect 490066 163898 497672 164134
rect 497908 163898 508278 164134
rect 508514 163898 516120 164134
rect 516356 163898 523962 164134
rect 524198 163898 531804 164134
rect 532040 163898 586302 164134
rect 586538 163898 586622 164134
rect 586858 163898 592650 164134
rect -8726 163866 592650 163898
rect -8726 158174 592650 158206
rect -8726 157938 -1974 158174
rect -1738 157938 -1654 158174
rect -1418 157938 48239 158174
rect 48475 157938 56081 158174
rect 56317 157938 63923 158174
rect 64159 157938 71765 158174
rect 72001 157938 82371 158174
rect 82607 157938 90213 158174
rect 90449 157938 98055 158174
rect 98291 157938 105897 158174
rect 106133 157938 149978 158174
rect 150214 157938 180698 158174
rect 180934 157938 277262 158174
rect 277498 157938 341539 158174
rect 341775 157938 349381 158174
rect 349617 157938 357223 158174
rect 357459 157938 365065 158174
rect 365301 157938 478067 158174
rect 478303 157938 485909 158174
rect 486145 157938 493751 158174
rect 493987 157938 501593 158174
rect 501829 157938 585342 158174
rect 585578 157938 585662 158174
rect 585898 157938 592650 158174
rect -8726 157854 592650 157938
rect -8726 157618 -1974 157854
rect -1738 157618 -1654 157854
rect -1418 157618 48239 157854
rect 48475 157618 56081 157854
rect 56317 157618 63923 157854
rect 64159 157618 71765 157854
rect 72001 157618 82371 157854
rect 82607 157618 90213 157854
rect 90449 157618 98055 157854
rect 98291 157618 105897 157854
rect 106133 157618 149978 157854
rect 150214 157618 180698 157854
rect 180934 157618 277262 157854
rect 277498 157618 341539 157854
rect 341775 157618 349381 157854
rect 349617 157618 357223 157854
rect 357459 157618 365065 157854
rect 365301 157618 478067 157854
rect 478303 157618 485909 157854
rect 486145 157618 493751 157854
rect 493987 157618 501593 157854
rect 501829 157618 585342 157854
rect 585578 157618 585662 157854
rect 585898 157618 592650 157854
rect -8726 157586 592650 157618
rect -8726 154454 592650 154486
rect -8726 154218 -2934 154454
rect -2698 154218 -2614 154454
rect -2378 154218 52160 154454
rect 52396 154218 60002 154454
rect 60238 154218 67844 154454
rect 68080 154218 75686 154454
rect 75922 154218 86292 154454
rect 86528 154218 94134 154454
rect 94370 154218 101976 154454
rect 102212 154218 109818 154454
rect 110054 154218 165338 154454
rect 165574 154218 277814 154454
rect 278050 154218 337618 154454
rect 337854 154218 345460 154454
rect 345696 154218 353302 154454
rect 353538 154218 361144 154454
rect 361380 154218 474146 154454
rect 474382 154218 481988 154454
rect 482224 154218 489830 154454
rect 490066 154218 497672 154454
rect 497908 154218 586302 154454
rect 586538 154218 586622 154454
rect 586858 154218 592650 154454
rect -8726 154134 592650 154218
rect -8726 153898 -2934 154134
rect -2698 153898 -2614 154134
rect -2378 153898 52160 154134
rect 52396 153898 60002 154134
rect 60238 153898 67844 154134
rect 68080 153898 75686 154134
rect 75922 153898 86292 154134
rect 86528 153898 94134 154134
rect 94370 153898 101976 154134
rect 102212 153898 109818 154134
rect 110054 153898 165338 154134
rect 165574 153898 277814 154134
rect 278050 153898 337618 154134
rect 337854 153898 345460 154134
rect 345696 153898 353302 154134
rect 353538 153898 361144 154134
rect 361380 153898 474146 154134
rect 474382 153898 481988 154134
rect 482224 153898 489830 154134
rect 490066 153898 497672 154134
rect 497908 153898 586302 154134
rect 586538 153898 586622 154134
rect 586858 153898 592650 154134
rect -8726 153866 592650 153898
rect -8726 148174 592650 148206
rect -8726 147938 -1974 148174
rect -1738 147938 -1654 148174
rect -1418 147938 48239 148174
rect 48475 147938 56081 148174
rect 56317 147938 63923 148174
rect 64159 147938 71765 148174
rect 72001 147938 82371 148174
rect 82607 147938 90213 148174
rect 90449 147938 98055 148174
rect 98291 147938 105897 148174
rect 106133 147938 149978 148174
rect 150214 147938 180698 148174
rect 180934 147938 277262 148174
rect 277498 147938 341539 148174
rect 341775 147938 349381 148174
rect 349617 147938 357223 148174
rect 357459 147938 365065 148174
rect 365301 147938 478067 148174
rect 478303 147938 485909 148174
rect 486145 147938 493751 148174
rect 493987 147938 501593 148174
rect 501829 147938 585342 148174
rect 585578 147938 585662 148174
rect 585898 147938 592650 148174
rect -8726 147854 592650 147938
rect -8726 147618 -1974 147854
rect -1738 147618 -1654 147854
rect -1418 147618 48239 147854
rect 48475 147618 56081 147854
rect 56317 147618 63923 147854
rect 64159 147618 71765 147854
rect 72001 147618 82371 147854
rect 82607 147618 90213 147854
rect 90449 147618 98055 147854
rect 98291 147618 105897 147854
rect 106133 147618 149978 147854
rect 150214 147618 180698 147854
rect 180934 147618 277262 147854
rect 277498 147618 341539 147854
rect 341775 147618 349381 147854
rect 349617 147618 357223 147854
rect 357459 147618 365065 147854
rect 365301 147618 478067 147854
rect 478303 147618 485909 147854
rect 486145 147618 493751 147854
rect 493987 147618 501593 147854
rect 501829 147618 585342 147854
rect 585578 147618 585662 147854
rect 585898 147618 592650 147854
rect -8726 147586 592650 147618
rect -8726 144454 592650 144486
rect -8726 144218 -2934 144454
rect -2698 144218 -2614 144454
rect -2378 144218 52160 144454
rect 52396 144218 60002 144454
rect 60238 144218 67844 144454
rect 68080 144218 75686 144454
rect 75922 144218 86292 144454
rect 86528 144218 94134 144454
rect 94370 144218 101976 144454
rect 102212 144218 109818 144454
rect 110054 144218 165338 144454
rect 165574 144218 277814 144454
rect 278050 144218 337618 144454
rect 337854 144218 345460 144454
rect 345696 144218 353302 144454
rect 353538 144218 361144 144454
rect 361380 144218 474146 144454
rect 474382 144218 481988 144454
rect 482224 144218 489830 144454
rect 490066 144218 497672 144454
rect 497908 144218 586302 144454
rect 586538 144218 586622 144454
rect 586858 144218 592650 144454
rect -8726 144134 592650 144218
rect -8726 143898 -2934 144134
rect -2698 143898 -2614 144134
rect -2378 143898 52160 144134
rect 52396 143898 60002 144134
rect 60238 143898 67844 144134
rect 68080 143898 75686 144134
rect 75922 143898 86292 144134
rect 86528 143898 94134 144134
rect 94370 143898 101976 144134
rect 102212 143898 109818 144134
rect 110054 143898 165338 144134
rect 165574 143898 277814 144134
rect 278050 143898 337618 144134
rect 337854 143898 345460 144134
rect 345696 143898 353302 144134
rect 353538 143898 361144 144134
rect 361380 143898 474146 144134
rect 474382 143898 481988 144134
rect 482224 143898 489830 144134
rect 490066 143898 497672 144134
rect 497908 143898 586302 144134
rect 586538 143898 586622 144134
rect 586858 143898 592650 144134
rect -8726 143866 592650 143898
rect -8726 138174 592650 138206
rect -8726 137938 -1974 138174
rect -1738 137938 -1654 138174
rect -1418 137938 48239 138174
rect 48475 137938 56081 138174
rect 56317 137938 63923 138174
rect 64159 137938 71765 138174
rect 72001 137938 82371 138174
rect 82607 137938 90213 138174
rect 90449 137938 98055 138174
rect 98291 137938 105897 138174
rect 106133 137938 149978 138174
rect 150214 137938 180698 138174
rect 180934 137938 211418 138174
rect 211654 137938 242138 138174
rect 242374 137938 272858 138174
rect 273094 137938 277262 138174
rect 277498 137938 341539 138174
rect 341775 137938 349381 138174
rect 349617 137938 357223 138174
rect 357459 137938 365065 138174
rect 365301 137938 478067 138174
rect 478303 137938 485909 138174
rect 486145 137938 493751 138174
rect 493987 137938 501593 138174
rect 501829 137938 585342 138174
rect 585578 137938 585662 138174
rect 585898 137938 592650 138174
rect -8726 137854 592650 137938
rect -8726 137618 -1974 137854
rect -1738 137618 -1654 137854
rect -1418 137618 48239 137854
rect 48475 137618 56081 137854
rect 56317 137618 63923 137854
rect 64159 137618 71765 137854
rect 72001 137618 82371 137854
rect 82607 137618 90213 137854
rect 90449 137618 98055 137854
rect 98291 137618 105897 137854
rect 106133 137618 149978 137854
rect 150214 137618 180698 137854
rect 180934 137618 211418 137854
rect 211654 137618 242138 137854
rect 242374 137618 272858 137854
rect 273094 137618 277262 137854
rect 277498 137618 341539 137854
rect 341775 137618 349381 137854
rect 349617 137618 357223 137854
rect 357459 137618 365065 137854
rect 365301 137618 478067 137854
rect 478303 137618 485909 137854
rect 486145 137618 493751 137854
rect 493987 137618 501593 137854
rect 501829 137618 585342 137854
rect 585578 137618 585662 137854
rect 585898 137618 592650 137854
rect -8726 137586 592650 137618
rect -8726 134454 592650 134486
rect -8726 134218 -2934 134454
rect -2698 134218 -2614 134454
rect -2378 134218 586302 134454
rect 586538 134218 586622 134454
rect 586858 134218 592650 134454
rect -8726 134134 592650 134218
rect -8726 133898 -2934 134134
rect -2698 133898 -2614 134134
rect -2378 133898 586302 134134
rect 586538 133898 586622 134134
rect 586858 133898 592650 134134
rect -8726 133866 592650 133898
rect -8726 128174 592650 128206
rect -8726 127938 -1974 128174
rect -1738 127938 -1654 128174
rect -1418 127938 13450 128174
rect 13686 127938 44170 128174
rect 44406 127938 74890 128174
rect 75126 127938 105610 128174
rect 105846 127938 136330 128174
rect 136566 127938 167050 128174
rect 167286 127938 197770 128174
rect 198006 127938 228490 128174
rect 228726 127938 259210 128174
rect 259446 127938 373098 128174
rect 373334 127938 403818 128174
rect 404054 127938 434538 128174
rect 434774 127938 448186 128174
rect 448422 127938 478906 128174
rect 479142 127938 509626 128174
rect 509862 127938 540346 128174
rect 540582 127938 571066 128174
rect 571302 127938 585342 128174
rect 585578 127938 585662 128174
rect 585898 127938 592650 128174
rect -8726 127854 592650 127938
rect -8726 127618 -1974 127854
rect -1738 127618 -1654 127854
rect -1418 127618 13450 127854
rect 13686 127618 44170 127854
rect 44406 127618 74890 127854
rect 75126 127618 105610 127854
rect 105846 127618 136330 127854
rect 136566 127618 167050 127854
rect 167286 127618 197770 127854
rect 198006 127618 228490 127854
rect 228726 127618 259210 127854
rect 259446 127618 373098 127854
rect 373334 127618 403818 127854
rect 404054 127618 434538 127854
rect 434774 127618 448186 127854
rect 448422 127618 478906 127854
rect 479142 127618 509626 127854
rect 509862 127618 540346 127854
rect 540582 127618 571066 127854
rect 571302 127618 585342 127854
rect 585578 127618 585662 127854
rect 585898 127618 592650 127854
rect -8726 127586 592650 127618
rect -8726 124454 592650 124486
rect -8726 124218 -2934 124454
rect -2698 124218 -2614 124454
rect -2378 124218 28810 124454
rect 29046 124218 59530 124454
rect 59766 124218 90250 124454
rect 90486 124218 120970 124454
rect 121206 124218 151690 124454
rect 151926 124218 182410 124454
rect 182646 124218 213130 124454
rect 213366 124218 243850 124454
rect 244086 124218 274570 124454
rect 274806 124218 388458 124454
rect 388694 124218 419178 124454
rect 419414 124218 463546 124454
rect 463782 124218 494266 124454
rect 494502 124218 524986 124454
rect 525222 124218 555706 124454
rect 555942 124218 586302 124454
rect 586538 124218 586622 124454
rect 586858 124218 592650 124454
rect -8726 124134 592650 124218
rect -8726 123898 -2934 124134
rect -2698 123898 -2614 124134
rect -2378 123898 28810 124134
rect 29046 123898 59530 124134
rect 59766 123898 90250 124134
rect 90486 123898 120970 124134
rect 121206 123898 151690 124134
rect 151926 123898 182410 124134
rect 182646 123898 213130 124134
rect 213366 123898 243850 124134
rect 244086 123898 274570 124134
rect 274806 123898 388458 124134
rect 388694 123898 419178 124134
rect 419414 123898 463546 124134
rect 463782 123898 494266 124134
rect 494502 123898 524986 124134
rect 525222 123898 555706 124134
rect 555942 123898 586302 124134
rect 586538 123898 586622 124134
rect 586858 123898 592650 124134
rect -8726 123866 592650 123898
rect -8726 118174 592650 118206
rect -8726 117938 -1974 118174
rect -1738 117938 -1654 118174
rect -1418 117938 13450 118174
rect 13686 117938 44170 118174
rect 44406 117938 74890 118174
rect 75126 117938 105610 118174
rect 105846 117938 136330 118174
rect 136566 117938 167050 118174
rect 167286 117938 197770 118174
rect 198006 117938 228490 118174
rect 228726 117938 259210 118174
rect 259446 117938 373098 118174
rect 373334 117938 403818 118174
rect 404054 117938 434538 118174
rect 434774 117938 448186 118174
rect 448422 117938 478906 118174
rect 479142 117938 509626 118174
rect 509862 117938 540346 118174
rect 540582 117938 571066 118174
rect 571302 117938 585342 118174
rect 585578 117938 585662 118174
rect 585898 117938 592650 118174
rect -8726 117854 592650 117938
rect -8726 117618 -1974 117854
rect -1738 117618 -1654 117854
rect -1418 117618 13450 117854
rect 13686 117618 44170 117854
rect 44406 117618 74890 117854
rect 75126 117618 105610 117854
rect 105846 117618 136330 117854
rect 136566 117618 167050 117854
rect 167286 117618 197770 117854
rect 198006 117618 228490 117854
rect 228726 117618 259210 117854
rect 259446 117618 373098 117854
rect 373334 117618 403818 117854
rect 404054 117618 434538 117854
rect 434774 117618 448186 117854
rect 448422 117618 478906 117854
rect 479142 117618 509626 117854
rect 509862 117618 540346 117854
rect 540582 117618 571066 117854
rect 571302 117618 585342 117854
rect 585578 117618 585662 117854
rect 585898 117618 592650 117854
rect -8726 117586 592650 117618
rect -8726 114454 592650 114486
rect -8726 114218 -2934 114454
rect -2698 114218 -2614 114454
rect -2378 114218 28810 114454
rect 29046 114218 59530 114454
rect 59766 114218 90250 114454
rect 90486 114218 120970 114454
rect 121206 114218 151690 114454
rect 151926 114218 182410 114454
rect 182646 114218 213130 114454
rect 213366 114218 243850 114454
rect 244086 114218 274570 114454
rect 274806 114218 388458 114454
rect 388694 114218 419178 114454
rect 419414 114218 463546 114454
rect 463782 114218 494266 114454
rect 494502 114218 524986 114454
rect 525222 114218 555706 114454
rect 555942 114218 586302 114454
rect 586538 114218 586622 114454
rect 586858 114218 592650 114454
rect -8726 114134 592650 114218
rect -8726 113898 -2934 114134
rect -2698 113898 -2614 114134
rect -2378 113898 28810 114134
rect 29046 113898 59530 114134
rect 59766 113898 90250 114134
rect 90486 113898 120970 114134
rect 121206 113898 151690 114134
rect 151926 113898 182410 114134
rect 182646 113898 213130 114134
rect 213366 113898 243850 114134
rect 244086 113898 274570 114134
rect 274806 113898 388458 114134
rect 388694 113898 419178 114134
rect 419414 113898 463546 114134
rect 463782 113898 494266 114134
rect 494502 113898 524986 114134
rect 525222 113898 555706 114134
rect 555942 113898 586302 114134
rect 586538 113898 586622 114134
rect 586858 113898 592650 114134
rect -8726 113866 592650 113898
rect -8726 108174 592650 108206
rect -8726 107938 -1974 108174
rect -1738 107938 -1654 108174
rect -1418 107938 13450 108174
rect 13686 107938 44170 108174
rect 44406 107938 74890 108174
rect 75126 107938 105610 108174
rect 105846 107938 136330 108174
rect 136566 107938 167050 108174
rect 167286 107938 197770 108174
rect 198006 107938 228490 108174
rect 228726 107938 259210 108174
rect 259446 107938 373098 108174
rect 373334 107938 403818 108174
rect 404054 107938 434538 108174
rect 434774 107938 448186 108174
rect 448422 107938 478906 108174
rect 479142 107938 509626 108174
rect 509862 107938 540346 108174
rect 540582 107938 571066 108174
rect 571302 107938 585342 108174
rect 585578 107938 585662 108174
rect 585898 107938 592650 108174
rect -8726 107854 592650 107938
rect -8726 107618 -1974 107854
rect -1738 107618 -1654 107854
rect -1418 107618 13450 107854
rect 13686 107618 44170 107854
rect 44406 107618 74890 107854
rect 75126 107618 105610 107854
rect 105846 107618 136330 107854
rect 136566 107618 167050 107854
rect 167286 107618 197770 107854
rect 198006 107618 228490 107854
rect 228726 107618 259210 107854
rect 259446 107618 373098 107854
rect 373334 107618 403818 107854
rect 404054 107618 434538 107854
rect 434774 107618 448186 107854
rect 448422 107618 478906 107854
rect 479142 107618 509626 107854
rect 509862 107618 540346 107854
rect 540582 107618 571066 107854
rect 571302 107618 585342 107854
rect 585578 107618 585662 107854
rect 585898 107618 592650 107854
rect -8726 107586 592650 107618
rect -8726 104454 592650 104486
rect -8726 104218 -2934 104454
rect -2698 104218 -2614 104454
rect -2378 104218 28810 104454
rect 29046 104218 59530 104454
rect 59766 104218 90250 104454
rect 90486 104218 120970 104454
rect 121206 104218 151690 104454
rect 151926 104218 182410 104454
rect 182646 104218 213130 104454
rect 213366 104218 243850 104454
rect 244086 104218 274570 104454
rect 274806 104218 388458 104454
rect 388694 104218 419178 104454
rect 419414 104218 463546 104454
rect 463782 104218 494266 104454
rect 494502 104218 524986 104454
rect 525222 104218 555706 104454
rect 555942 104218 586302 104454
rect 586538 104218 586622 104454
rect 586858 104218 592650 104454
rect -8726 104134 592650 104218
rect -8726 103898 -2934 104134
rect -2698 103898 -2614 104134
rect -2378 103898 28810 104134
rect 29046 103898 59530 104134
rect 59766 103898 90250 104134
rect 90486 103898 120970 104134
rect 121206 103898 151690 104134
rect 151926 103898 182410 104134
rect 182646 103898 213130 104134
rect 213366 103898 243850 104134
rect 244086 103898 274570 104134
rect 274806 103898 388458 104134
rect 388694 103898 419178 104134
rect 419414 103898 463546 104134
rect 463782 103898 494266 104134
rect 494502 103898 524986 104134
rect 525222 103898 555706 104134
rect 555942 103898 586302 104134
rect 586538 103898 586622 104134
rect 586858 103898 592650 104134
rect -8726 103866 592650 103898
rect -8726 98174 592650 98206
rect -8726 97938 -1974 98174
rect -1738 97938 -1654 98174
rect -1418 97938 13450 98174
rect 13686 97938 44170 98174
rect 44406 97938 74890 98174
rect 75126 97938 105610 98174
rect 105846 97938 136330 98174
rect 136566 97938 167050 98174
rect 167286 97938 197770 98174
rect 198006 97938 228490 98174
rect 228726 97938 259210 98174
rect 259446 97938 373098 98174
rect 373334 97938 403818 98174
rect 404054 97938 434538 98174
rect 434774 97938 448186 98174
rect 448422 97938 478906 98174
rect 479142 97938 509626 98174
rect 509862 97938 540346 98174
rect 540582 97938 571066 98174
rect 571302 97938 585342 98174
rect 585578 97938 585662 98174
rect 585898 97938 592650 98174
rect -8726 97854 592650 97938
rect -8726 97618 -1974 97854
rect -1738 97618 -1654 97854
rect -1418 97618 13450 97854
rect 13686 97618 44170 97854
rect 44406 97618 74890 97854
rect 75126 97618 105610 97854
rect 105846 97618 136330 97854
rect 136566 97618 167050 97854
rect 167286 97618 197770 97854
rect 198006 97618 228490 97854
rect 228726 97618 259210 97854
rect 259446 97618 373098 97854
rect 373334 97618 403818 97854
rect 404054 97618 434538 97854
rect 434774 97618 448186 97854
rect 448422 97618 478906 97854
rect 479142 97618 509626 97854
rect 509862 97618 540346 97854
rect 540582 97618 571066 97854
rect 571302 97618 585342 97854
rect 585578 97618 585662 97854
rect 585898 97618 592650 97854
rect -8726 97586 592650 97618
rect -8726 94454 592650 94486
rect -8726 94218 -2934 94454
rect -2698 94218 -2614 94454
rect -2378 94218 28810 94454
rect 29046 94218 59530 94454
rect 59766 94218 90250 94454
rect 90486 94218 120970 94454
rect 121206 94218 151690 94454
rect 151926 94218 182410 94454
rect 182646 94218 213130 94454
rect 213366 94218 243850 94454
rect 244086 94218 274570 94454
rect 274806 94218 388458 94454
rect 388694 94218 419178 94454
rect 419414 94218 463546 94454
rect 463782 94218 494266 94454
rect 494502 94218 524986 94454
rect 525222 94218 555706 94454
rect 555942 94218 586302 94454
rect 586538 94218 586622 94454
rect 586858 94218 592650 94454
rect -8726 94134 592650 94218
rect -8726 93898 -2934 94134
rect -2698 93898 -2614 94134
rect -2378 93898 28810 94134
rect 29046 93898 59530 94134
rect 59766 93898 90250 94134
rect 90486 93898 120970 94134
rect 121206 93898 151690 94134
rect 151926 93898 182410 94134
rect 182646 93898 213130 94134
rect 213366 93898 243850 94134
rect 244086 93898 274570 94134
rect 274806 93898 388458 94134
rect 388694 93898 419178 94134
rect 419414 93898 463546 94134
rect 463782 93898 494266 94134
rect 494502 93898 524986 94134
rect 525222 93898 555706 94134
rect 555942 93898 586302 94134
rect 586538 93898 586622 94134
rect 586858 93898 592650 94134
rect -8726 93866 592650 93898
rect -8726 88174 592650 88206
rect -8726 87938 -1974 88174
rect -1738 87938 -1654 88174
rect -1418 87938 585342 88174
rect 585578 87938 585662 88174
rect 585898 87938 592650 88174
rect -8726 87854 592650 87938
rect -8726 87618 -1974 87854
rect -1738 87618 -1654 87854
rect -1418 87618 585342 87854
rect 585578 87618 585662 87854
rect 585898 87618 592650 87854
rect -8726 87586 592650 87618
rect -8726 84454 592650 84486
rect -8726 84218 -2934 84454
rect -2698 84218 -2614 84454
rect -2378 84218 586302 84454
rect 586538 84218 586622 84454
rect 586858 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -2934 84134
rect -2698 83898 -2614 84134
rect -2378 83898 586302 84134
rect 586538 83898 586622 84134
rect 586858 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 78174 592650 78206
rect -8726 77938 -1974 78174
rect -1738 77938 -1654 78174
rect -1418 77938 585342 78174
rect 585578 77938 585662 78174
rect 585898 77938 592650 78174
rect -8726 77854 592650 77938
rect -8726 77618 -1974 77854
rect -1738 77618 -1654 77854
rect -1418 77618 585342 77854
rect 585578 77618 585662 77854
rect 585898 77618 592650 77854
rect -8726 77586 592650 77618
rect -8726 74454 592650 74486
rect -8726 74218 -2934 74454
rect -2698 74218 -2614 74454
rect -2378 74218 586302 74454
rect 586538 74218 586622 74454
rect 586858 74218 592650 74454
rect -8726 74134 592650 74218
rect -8726 73898 -2934 74134
rect -2698 73898 -2614 74134
rect -2378 73898 586302 74134
rect 586538 73898 586622 74134
rect 586858 73898 592650 74134
rect -8726 73866 592650 73898
rect -8726 68174 592650 68206
rect -8726 67938 -1974 68174
rect -1738 67938 -1654 68174
rect -1418 67938 585342 68174
rect 585578 67938 585662 68174
rect 585898 67938 592650 68174
rect -8726 67854 592650 67938
rect -8726 67618 -1974 67854
rect -1738 67618 -1654 67854
rect -1418 67618 585342 67854
rect 585578 67618 585662 67854
rect 585898 67618 592650 67854
rect -8726 67586 592650 67618
rect -8726 64454 592650 64486
rect -8726 64218 -2934 64454
rect -2698 64218 -2614 64454
rect -2378 64218 586302 64454
rect 586538 64218 586622 64454
rect 586858 64218 592650 64454
rect -8726 64171 592650 64218
rect -8726 64134 293034 64171
rect -8726 63898 -2934 64134
rect -2698 63898 -2614 64134
rect -2378 63935 293034 64134
rect 293270 64134 592650 64171
rect 293270 63935 586302 64134
rect -2378 63898 586302 63935
rect 586538 63898 586622 64134
rect 586858 63898 592650 64134
rect -8726 63866 592650 63898
rect -8726 58174 592650 58206
rect -8726 57938 -1974 58174
rect -1738 57938 -1654 58174
rect -1418 57938 277674 58174
rect 277910 57938 308394 58174
rect 308630 57938 585342 58174
rect 585578 57938 585662 58174
rect 585898 57938 592650 58174
rect -8726 57854 592650 57938
rect -8726 57618 -1974 57854
rect -1738 57618 -1654 57854
rect -1418 57618 277674 57854
rect 277910 57618 308394 57854
rect 308630 57618 585342 57854
rect 585578 57618 585662 57854
rect 585898 57618 592650 57854
rect -8726 57586 592650 57618
rect -8726 54454 592650 54486
rect -8726 54218 -2934 54454
rect -2698 54218 -2614 54454
rect -2378 54218 293034 54454
rect 293270 54218 586302 54454
rect 586538 54218 586622 54454
rect 586858 54218 592650 54454
rect -8726 54134 592650 54218
rect -8726 53898 -2934 54134
rect -2698 53898 -2614 54134
rect -2378 53898 293034 54134
rect 293270 53898 586302 54134
rect 586538 53898 586622 54134
rect 586858 53898 592650 54134
rect -8726 53866 592650 53898
rect -8726 48174 592650 48206
rect -8726 47938 -1974 48174
rect -1738 47938 -1654 48174
rect -1418 47938 277674 48174
rect 277910 47938 308394 48174
rect 308630 47938 585342 48174
rect 585578 47938 585662 48174
rect 585898 47938 592650 48174
rect -8726 47854 592650 47938
rect -8726 47618 -1974 47854
rect -1738 47618 -1654 47854
rect -1418 47618 277674 47854
rect 277910 47618 308394 47854
rect 308630 47618 585342 47854
rect 585578 47618 585662 47854
rect 585898 47618 592650 47854
rect -8726 47586 592650 47618
rect -8726 44454 592650 44486
rect -8726 44218 -2934 44454
rect -2698 44218 -2614 44454
rect -2378 44218 293034 44454
rect 293270 44218 586302 44454
rect 586538 44218 586622 44454
rect 586858 44218 592650 44454
rect -8726 44134 592650 44218
rect -8726 43898 -2934 44134
rect -2698 43898 -2614 44134
rect -2378 43898 293034 44134
rect 293270 43898 586302 44134
rect 586538 43898 586622 44134
rect 586858 43898 592650 44134
rect -8726 43866 592650 43898
rect -8726 38174 592650 38206
rect -8726 37938 -1974 38174
rect -1738 37938 -1654 38174
rect -1418 37938 277674 38174
rect 277910 37938 308394 38174
rect 308630 37938 585342 38174
rect 585578 37938 585662 38174
rect 585898 37938 592650 38174
rect -8726 37854 592650 37938
rect -8726 37618 -1974 37854
rect -1738 37618 -1654 37854
rect -1418 37618 277674 37854
rect 277910 37618 308394 37854
rect 308630 37618 585342 37854
rect 585578 37618 585662 37854
rect 585898 37618 592650 37854
rect -8726 37586 592650 37618
rect -8726 34454 592650 34486
rect -8726 34218 -2934 34454
rect -2698 34218 -2614 34454
rect -2378 34218 293034 34454
rect 293270 34218 586302 34454
rect 586538 34218 586622 34454
rect 586858 34218 592650 34454
rect -8726 34134 592650 34218
rect -8726 33898 -2934 34134
rect -2698 33898 -2614 34134
rect -2378 33898 293034 34134
rect 293270 33898 586302 34134
rect 586538 33898 586622 34134
rect 586858 33898 592650 34134
rect -8726 33866 592650 33898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use tt_um_as1802  tt_top1.branch\[0\].col_um\[0\].um_bot_I.block_0_0.tt_um_I
timestamp 0
transform 1 0 9200 0 1 90848
box 1066 2 271438 44064
use tt_um_loopback  tt_top1.branch\[0\].col_um\[0\].um_top_I.block_1_0.tt_um_I
timestamp 0
transform 1 0 9200 0 -1 212704
box 1066 1040 32632 21760
use tt_um_urish_simon  tt_top1.branch\[0\].col_um\[1\].um_bot_I.block_0_1.tt_um_I
timestamp 0
transform 1 0 43332 0 1 134912
box 1066 1040 32632 44064
use tt_um_power_test  tt_top1.branch\[0\].col_um\[1\].um_top_I.block_1_1.tt_um_I
timestamp 0
transform 1 0 43332 0 -1 212704
box -1084 -6172 32992 21760
use tt_um_kiwih_tt_top  tt_top1.branch\[0\].col_um\[2\].um_bot_I.block_0_2.tt_um_I
timestamp 0
transform 1 0 77464 0 1 134912
box 1066 1040 32632 44064
use tt_um_htfab_totp  tt_top1.branch\[0\].col_um\[2\].um_top_I.block_1_2.tt_um_I
timestamp 0
transform 1 0 77464 0 -1 279072
box 106 2 67698 44064
use tt_um_wokwi_366318576852367361  tt_top1.branch\[0\].col_um\[3\].um_bot_I.block_0_3.tt_um_I
timestamp 0
transform 1 0 111596 0 1 157216
box 1066 1040 32632 21760
use tt_um_gatecat_fpga_top  tt_top1.branch\[0\].col_um\[3\].um_top_I.block_1_3.tt_um_I
timestamp 0
transform 1 0 111596 0 -1 235008
box 1066 1040 32830 44064
use tt_um_urish_dffram  tt_top1.branch\[0\].col_um\[4\].um_bot_I.block_0_4.tt_um_I
timestamp 0
transform 1 0 145728 0 1 134912
box 1066 1040 134910 44064
use tt_um_Reloj_top  tt_top1.branch\[0\].col_um\[4\].um_top_I.block_1_4.tt_um_I
timestamp 0
transform 1 0 145728 0 -1 279072
box 1066 1040 66646 44064
use tt_um_algofoogle_solo_squash  tt_top1.branch\[0\].col_um\[5\].um_top_I.block_1_5.tt_um_I
timestamp 0
transform 1 0 179860 0 -1 212704
box 1066 1040 32632 21760
use tt_um_apu_pulse  tt_top1.branch\[0\].col_um\[6\].um_top_I.block_1_6.tt_um_I
timestamp 0
transform 1 0 213992 0 -1 212704
box 13 274 33566 21760
use tt_um_thorkn_vgaclock  tt_top1.branch\[0\].col_um\[7\].um_top_I.block_1_7.tt_um_I
timestamp 0
transform 1 0 248124 0 -1 212704
box 1066 1040 32632 21760
use tt_mux  tt_top1.branch\[0\].mux_I
timestamp 0
transform 1 0 9200 0 1 179520
box 750 0 272504 10880
use tt_um_greycode_top  tt_top1.branch\[1\].col_um\[0\].um_bot_I.block_0_16.tt_um_I
timestamp 0
transform -1 0 575552 0 1 90848
box 1066 1040 134910 44064
use tt_um_loopback  tt_top1.branch\[1\].col_um\[0\].um_top_I.block_1_16.tt_um_I
timestamp 0
transform -1 0 575000 0 -1 212704
box 1066 1040 32632 21760
use tt_um_moyes0_top_module  tt_top1.branch\[1\].col_um\[1\].um_bot_I.block_0_17.tt_um_I
timestamp 0
transform -1 0 540868 0 1 157216
box 1066 1040 32632 21760
use tt_um_wokwi_347497504164545108  tt_top1.branch\[1\].col_um\[1\].um_top_I.block_1_17.tt_um_I
timestamp 0
transform -1 0 540868 0 -1 212704
box 1066 1040 32632 21760
use tt_um_vga_clock  tt_top1.branch\[1\].col_um\[2\].um_bot_I.block_0_18.tt_um_I
timestamp 0
transform -1 0 506736 0 1 134912
box 1066 1040 32632 44064
use tt_um_wokwi_347144898258928211  tt_top1.branch\[1\].col_um\[2\].um_top_I.block_1_18.tt_um_I
timestamp 0
transform -1 0 506736 0 -1 212704
box 1066 1040 32632 21760
use tt_um_TrainLED2_top  tt_top1.branch\[1\].col_um\[3\].um_bot_I.block_0_19.tt_um_I
timestamp 0
transform -1 0 472604 0 1 157216
box 1066 1040 32632 21760
use tt_um_wokwi_347417602591556180  tt_top1.branch\[1\].col_um\[3\].um_top_I.block_1_19.tt_um_I
timestamp 0
transform -1 0 472604 0 -1 212704
box 1066 1040 32632 21760
use tt_um_tomkeddie_a  tt_top1.branch\[1\].col_um\[4\].um_bot_I.block_0_20.tt_um_I
timestamp 0
transform -1 0 439024 0 1 90848
box 1066 1040 66646 44064
use tt_um_millerresearch_top  tt_top1.branch\[1\].col_um\[4\].um_top_I.block_1_20.tt_um_I
timestamp 0
transform -1 0 438472 0 -1 235008
box 1066 1040 32632 44064
use tt_um_ternaryPC_radixconvert  tt_top1.branch\[1\].col_um\[5\].um_bot_I.block_0_21.tt_um_I
timestamp 0
transform -1 0 404340 0 1 157216
box 1066 1040 32632 21760
use tt_um_psychogenic_neptuneproportional  tt_top1.branch\[1\].col_um\[5\].um_top_I.block_1_21.tt_um_I
timestamp 0
transform -1 0 404340 0 -1 212704
box 1066 1040 32632 21760
use tt_um_MichaelBell_hovalaag  tt_top1.branch\[1\].col_um\[6\].um_bot_I.block_0_22.tt_um_I
timestamp 0
transform -1 0 370208 0 1 134912
box 1066 1040 32632 44064
use tt_um_test  tt_top1.branch\[1\].col_um\[6\].um_top_I.block_1_22.tt_um_I
timestamp 0
transform -1 0 370208 0 -1 212704
box 1066 1040 32632 21760
use tt_um_cam  tt_top1.branch\[1\].col_um\[7\].um_bot_I.block_0_23.tt_um_I
timestamp 0
transform -1 0 336076 0 1 157216
box 1066 1040 32632 21760
use sky130_sram_2kbyte_1rw1r_32x512_8  tt_top1.branch\[1\].col_um\[7\].um_top_I.block_1_23.sram
timestamp 0
transform 1 0 302496 0 1 240000
box 0 0 136620 83308
use tt_um_urish_sram_poc  tt_top1.branch\[1\].col_um\[7\].um_top_I.block_1_23.tt_um_I
timestamp 0
transform -1 0 336076 0 -1 212704
box 1066 0 32632 21760
use tt_mux  tt_top1.branch\[1\].mux_I
timestamp 0
transform -1 0 575000 0 1 179520
box 750 0 272504 10880
use tt_ctrl  tt_top1.ctrl_I
timestamp 0
transform 1 0 273424 0 1 21760
box 790 0 36010 44064
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 37586 592650 38206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 47586 592650 48206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 57586 592650 58206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 67586 592650 68206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 77586 592650 78206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 87586 592650 88206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 97586 592650 98206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 107586 592650 108206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 117586 592650 118206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 127586 592650 128206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 137586 592650 138206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 147586 592650 148206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 157586 592650 158206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 167586 592650 168206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 177586 592650 178206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 187586 592650 188206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 197586 592650 198206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 207586 592650 208206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 217586 592650 218206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 227586 592650 228206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 237586 592650 238206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 247586 592650 248206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 257586 592650 258206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 267586 592650 268206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 277586 592650 278206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 287586 592650 288206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 297586 592650 298206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 307586 592650 308206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 317586 592650 318206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 327586 592650 328206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 337586 592650 338206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 347586 592650 348206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 357586 592650 358206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 367586 592650 368206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 377586 592650 378206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 387586 592650 388206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 397586 592650 398206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 407586 592650 408206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 417586 592650 418206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 427586 592650 428206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 437586 592650 438206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 447586 592650 448206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 457586 592650 458206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 467586 592650 468206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 477586 592650 478206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 487586 592650 488206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 497586 592650 498206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 507586 592650 508206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 517586 592650 518206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 527586 592650 528206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 537586 592650 538206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 547586 592650 548206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 557586 592650 558206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 567586 592650 568206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 577586 592650 578206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 587586 592650 588206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 597586 592650 598206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 607586 592650 608206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 617586 592650 618206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 627586 592650 628206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 637586 592650 638206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 647586 592650 648206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 657586 592650 658206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 667586 592650 668206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 677586 592650 678206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 687586 592650 688206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 697586 592650 698206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 33866 592650 34486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43866 592650 44486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 53866 592650 54486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 63866 592650 64486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 73866 592650 74486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 93866 592650 94486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 103866 592650 104486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 113866 592650 114486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 123866 592650 124486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 133866 592650 134486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 143866 592650 144486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 153866 592650 154486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 163866 592650 164486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 183866 592650 184486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 193866 592650 194486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 203866 592650 204486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 213866 592650 214486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223866 592650 224486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 233866 592650 234486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 243866 592650 244486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 253866 592650 254486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 273866 592650 274486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 283866 592650 284486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 293866 592650 294486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 303866 592650 304486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 313866 592650 314486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 323866 592650 324486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 333866 592650 334486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 343866 592650 344486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 363866 592650 364486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 373866 592650 374486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 383866 592650 384486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 393866 592650 394486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403866 592650 404486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 413866 592650 414486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 423866 592650 424486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 433866 592650 434486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 453866 592650 454486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 463866 592650 464486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 473866 592650 474486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 483866 592650 484486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 493866 592650 494486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 503866 592650 504486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 513866 592650 514486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 523866 592650 524486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 543866 592650 544486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 553866 592650 554486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 563866 592650 564486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 573866 592650 574486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583866 592650 584486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 593866 592650 594486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 603866 592650 604486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 613866 592650 614486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 633866 592650 634486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 643866 592650 644486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 653866 592650 654486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 663866 592650 664486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 673866 592650 674486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 683866 592650 684486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 693866 592650 694486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
